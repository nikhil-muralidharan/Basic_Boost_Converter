magic
tech sky130A
timestamp 1660758149
<< nwell >>
rect -205 115 405 280
<< pmoslvt >>
rect -55 145 -20 245
rect 30 145 65 245
rect 215 145 250 245
<< nmoslvt >>
rect -55 -325 -40 -225
rect 90 -325 105 -225
rect 235 -325 250 -225
<< ndiff >>
rect -105 -240 -55 -225
rect -105 -310 -90 -240
rect -70 -310 -55 -240
rect -105 -325 -55 -310
rect -40 -240 10 -225
rect -40 -310 -25 -240
rect -5 -310 10 -240
rect -40 -325 10 -310
rect 40 -240 90 -225
rect 40 -310 55 -240
rect 75 -310 90 -240
rect 40 -325 90 -310
rect 105 -240 155 -225
rect 105 -310 120 -240
rect 140 -310 155 -240
rect 105 -325 155 -310
rect 185 -240 235 -225
rect 185 -310 200 -240
rect 220 -310 235 -240
rect 185 -325 235 -310
rect 250 -240 300 -225
rect 250 -310 265 -240
rect 285 -310 300 -240
rect 250 -325 300 -310
<< pdiff >>
rect -105 230 -55 245
rect -105 160 -90 230
rect -70 160 -55 230
rect -105 145 -55 160
rect -20 230 30 245
rect -20 160 -5 230
rect 15 160 30 230
rect -20 145 30 160
rect 65 230 115 245
rect 65 160 80 230
rect 100 160 115 230
rect 65 145 115 160
rect 165 230 215 245
rect 165 160 180 230
rect 200 160 215 230
rect 165 145 215 160
rect 250 230 300 245
rect 250 160 265 230
rect 285 160 300 230
rect 250 145 300 160
<< ndiffc >>
rect -90 -310 -70 -240
rect -25 -310 -5 -240
rect 55 -310 75 -240
rect 120 -310 140 -240
rect 200 -310 220 -240
rect 265 -310 285 -240
<< pdiffc >>
rect -90 160 -70 230
rect -5 160 15 230
rect 80 160 100 230
rect 180 160 200 230
rect 265 160 285 230
<< psubdiff >>
rect -185 -240 -135 -225
rect -185 -310 -170 -240
rect -150 -310 -135 -240
rect -185 -325 -135 -310
<< nsubdiff >>
rect -185 230 -135 245
rect -185 160 -170 230
rect -150 160 -135 230
rect -185 145 -135 160
<< psubdiffcont >>
rect -170 -310 -150 -240
<< nsubdiffcont >>
rect -170 160 -150 230
<< poly >>
rect -55 245 -20 260
rect 30 245 65 260
rect 215 245 250 260
rect -55 130 -20 145
rect 30 130 65 145
rect 215 130 250 145
rect -55 115 -40 130
rect -80 105 -40 115
rect -80 85 -70 105
rect -50 85 -40 105
rect -80 75 -40 85
rect 50 55 65 130
rect 210 120 250 130
rect 210 100 220 120
rect 240 100 250 120
rect 210 90 250 100
rect 50 45 90 55
rect 50 25 60 45
rect 80 25 90 45
rect 50 15 90 25
rect -80 -180 -40 -170
rect -80 -200 -70 -180
rect -50 -200 -40 -180
rect -80 -210 -40 -200
rect 65 -180 105 -170
rect 65 -200 75 -180
rect 95 -200 105 -180
rect 65 -210 105 -200
rect 210 -180 250 -170
rect 210 -200 220 -180
rect 240 -200 250 -180
rect 210 -210 250 -200
rect -55 -225 -40 -210
rect 90 -225 105 -210
rect 235 -225 250 -210
rect -55 -340 -40 -325
rect 90 -340 105 -325
rect 235 -340 250 -325
rect -55 -350 -15 -340
rect -55 -370 -45 -350
rect -25 -370 -15 -350
rect -55 -380 -15 -370
rect 90 -350 130 -340
rect 90 -370 100 -350
rect 120 -370 130 -350
rect 90 -380 130 -370
<< polycont >>
rect -70 85 -50 105
rect 220 100 240 120
rect 60 25 80 45
rect -70 -200 -50 -180
rect 75 -200 95 -180
rect 220 -200 240 -180
rect -45 -370 -25 -350
rect 100 -370 120 -350
<< locali >>
rect -180 230 -140 240
rect -180 160 -170 230
rect -150 160 -140 230
rect -180 150 -140 160
rect -100 230 -60 240
rect -100 160 -90 230
rect -70 160 -60 230
rect -100 150 -60 160
rect -15 230 25 240
rect -15 160 -5 230
rect 15 160 25 230
rect -15 150 25 160
rect 70 230 110 240
rect 70 160 80 230
rect 100 160 110 230
rect 70 150 110 160
rect 170 230 210 240
rect 170 160 180 230
rect 200 160 210 230
rect 170 150 210 160
rect 255 230 295 240
rect 255 160 265 230
rect 285 160 295 230
rect 255 150 295 160
rect -80 105 -40 115
rect -80 85 -70 105
rect -50 85 -40 105
rect 80 95 100 150
rect 210 120 250 130
rect 210 100 220 120
rect 240 100 250 120
rect 210 95 250 100
rect -80 75 -40 85
rect -15 75 250 95
rect 275 100 295 150
rect 275 80 375 100
rect -70 -170 -50 75
rect -80 -180 -40 -170
rect -80 -200 -70 -180
rect -50 -200 -40 -180
rect -80 -210 -40 -200
rect -15 -230 5 75
rect 50 45 90 55
rect 50 25 60 45
rect 80 25 90 45
rect 50 15 90 25
rect 65 -170 90 15
rect 65 -180 105 -170
rect 65 -200 75 -180
rect 95 -200 105 -180
rect 65 -210 105 -200
rect 130 -230 150 75
rect 220 -170 240 75
rect 210 -180 250 -170
rect 210 -200 220 -180
rect 240 -200 250 -180
rect 210 -210 250 -200
rect 275 -230 295 80
rect -180 -240 -140 -230
rect -180 -310 -170 -240
rect -150 -310 -140 -240
rect -180 -320 -140 -310
rect -100 -240 -60 -230
rect -100 -310 -90 -240
rect -70 -310 -60 -240
rect -100 -320 -60 -310
rect -35 -240 5 -230
rect -35 -310 -25 -240
rect -5 -310 5 -240
rect -35 -320 5 -310
rect 45 -240 85 -230
rect 45 -310 55 -240
rect 75 -310 85 -240
rect 45 -320 85 -310
rect 110 -240 150 -230
rect 110 -310 120 -240
rect 140 -310 150 -240
rect 110 -320 150 -310
rect 190 -240 230 -230
rect 190 -310 200 -240
rect 220 -310 230 -240
rect 190 -320 230 -310
rect 255 -240 295 -230
rect 255 -310 265 -240
rect 285 -310 295 -240
rect 255 -320 295 -310
rect 355 -340 375 80
rect -55 -350 -15 -340
rect -55 -370 -45 -350
rect -25 -370 -15 -350
rect -55 -380 -15 -370
rect 90 -350 130 -340
rect 90 -370 100 -350
rect 120 -370 130 -350
rect 355 -360 410 -340
rect 90 -380 130 -370
<< viali >>
rect -170 160 -150 230
rect -90 160 -70 230
rect 180 160 200 230
rect -170 -310 -150 -240
rect -90 -310 -70 -240
rect 55 -310 75 -240
rect 200 -310 220 -240
<< metal1 >>
rect -205 230 405 240
rect -205 160 -170 230
rect -150 160 -90 230
rect -70 160 180 230
rect 200 160 405 230
rect -205 150 405 160
rect -205 -240 405 -230
rect -205 -310 -170 -240
rect -150 -310 -90 -240
rect -70 -310 55 -240
rect 75 -310 200 -240
rect 220 -310 405 -240
rect -205 -320 405 -310
<< labels >>
rlabel metal1 -205 195 -205 195 7 VP
port 1 w
rlabel locali 335 90 335 90 3 Y
port 5 e
rlabel metal1 -205 -275 -205 -275 7 VN
port 2 w
rlabel locali -35 -380 -35 -380 5 A
port 3 s
rlabel locali 110 -380 110 -380 5 B
port 4 s
<< end >>
