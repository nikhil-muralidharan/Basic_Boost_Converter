magic
tech sky130A
timestamp 1658392951
<< nwell >>
rect -618 219 -179 246
rect -620 96 -179 219
rect -455 95 -179 96
<< pmoslvt >>
rect -455 125 -420 220
rect -290 125 -255 220
<< nmoslvt >>
rect -440 -80 -425 15
rect -375 -80 -359 15
<< ndiff >>
rect -492 -5 -440 15
rect -492 -61 -475 -5
rect -454 -61 -440 -5
rect -492 -80 -440 -61
rect -425 -5 -375 15
rect -425 -61 -410 -5
rect -389 -61 -375 -5
rect -425 -80 -375 -61
rect -359 -5 -304 15
rect -359 -61 -340 -5
rect -319 -61 -304 -5
rect -359 -80 -304 -61
<< pdiff >>
rect -505 219 -455 220
rect -506 200 -455 219
rect -506 145 -489 200
rect -468 145 -455 200
rect -506 125 -455 145
rect -420 219 -370 220
rect -420 199 -369 219
rect -420 144 -405 199
rect -384 144 -369 199
rect -420 125 -369 144
rect -342 200 -290 220
rect -342 145 -325 200
rect -304 145 -290 200
rect -342 125 -290 145
rect -255 201 -200 220
rect -255 145 -235 201
rect -214 145 -200 201
rect -255 125 -200 145
<< ndiffc >>
rect -475 -61 -454 -5
rect -410 -61 -389 -5
rect -340 -61 -319 -5
<< pdiffc >>
rect -489 145 -468 200
rect -405 144 -384 199
rect -325 145 -304 200
rect -235 145 -214 201
<< psubdiff >>
rect -571 -5 -519 15
rect -571 -61 -555 -5
rect -534 -61 -519 -5
rect -571 -80 -519 -61
<< nsubdiff >>
rect -596 200 -545 220
rect -596 145 -581 200
rect -560 145 -545 200
rect -596 125 -545 145
<< psubdiffcont >>
rect -555 -61 -534 -5
<< nsubdiffcont >>
rect -581 145 -560 200
<< poly >>
rect -455 220 -420 246
rect -290 220 -255 245
rect -455 95 -420 125
rect -290 95 -255 125
rect -455 70 -439 95
rect -395 70 -359 75
rect -285 70 -270 95
rect -455 55 -425 70
rect -440 15 -425 55
rect -395 68 -270 70
rect -395 48 -387 68
rect -368 55 -270 68
rect -368 48 -359 55
rect -395 40 -359 48
rect -375 15 -359 40
rect -440 -95 -425 -80
rect -375 -95 -359 -80
rect -465 -102 -425 -95
rect -465 -122 -455 -102
rect -436 -122 -425 -102
rect -465 -130 -425 -122
<< polycont >>
rect -387 48 -368 68
rect -455 -122 -436 -102
<< locali >>
rect -590 200 -551 215
rect -590 145 -581 200
rect -560 145 -551 200
rect -590 130 -551 145
rect -499 200 -460 215
rect -499 145 -489 200
rect -468 145 -460 200
rect -499 130 -460 145
rect -415 199 -376 215
rect -415 144 -405 199
rect -384 144 -376 199
rect -415 130 -376 144
rect -335 200 -295 215
rect -335 145 -325 200
rect -304 145 -295 200
rect -335 130 -295 145
rect -245 201 -205 215
rect -245 145 -235 201
rect -214 145 -205 201
rect -245 130 -205 145
rect -480 65 -460 130
rect -395 68 -359 75
rect -395 65 -387 68
rect -480 48 -387 65
rect -368 48 -359 68
rect -235 65 -215 130
rect -260 50 -179 65
rect -480 45 -359 48
rect -480 10 -460 45
rect -395 40 -359 45
rect -335 45 -179 50
rect -335 30 -240 45
rect -335 10 -315 30
rect -565 -5 -525 10
rect -565 -61 -555 -5
rect -534 -61 -525 -5
rect -565 -75 -525 -61
rect -485 -5 -445 10
rect -485 -61 -475 -5
rect -454 -61 -445 -5
rect -485 -75 -445 -61
rect -420 -5 -380 10
rect -335 9 -310 10
rect -420 -61 -410 -5
rect -389 -61 -380 -5
rect -420 -75 -380 -61
rect -350 -5 -310 9
rect -350 -61 -340 -5
rect -319 -61 -310 -5
rect -350 -75 -310 -61
rect -465 -100 -425 -95
rect -620 -102 -425 -100
rect -620 -120 -455 -102
rect -465 -122 -455 -120
rect -436 -122 -425 -102
rect -465 -130 -425 -122
<< viali >>
rect -405 144 -384 199
rect -325 145 -304 200
rect -555 -61 -534 -5
rect -340 -61 -319 -5
<< metal1 >>
rect -620 200 -180 215
rect -620 199 -325 200
rect -620 144 -405 199
rect -384 145 -325 199
rect -304 145 -180 200
rect -384 144 -180 145
rect -620 130 -180 144
rect -620 -5 -310 10
rect -620 -61 -555 -5
rect -534 -61 -340 -5
rect -319 -61 -310 -5
rect -620 -75 -310 -61
rect -304 -75 -179 10
<< rmetal1 >>
rect -310 -75 -304 10
<< labels >>
rlabel metal1 -620 170 -620 170 7 Vdd
port 3 w
rlabel metal1 -620 -35 -620 -35 7 Gnd
port 4 w
rlabel locali -620 -110 -620 -110 7 in
port 1 w
rlabel locali -179 55 -179 55 3 out
port 2 e
<< end >>
