magic
tech sky130A
timestamp 1659595967
<< nwell >>
rect -140 -50 470 175
<< pmoslvt >>
rect 30 5 65 105
rect 115 5 150 105
rect 280 5 315 105
<< nmoslvt >>
rect 30 -280 45 -180
rect 95 -280 110 -180
rect 280 -280 295 -180
rect 345 -280 360 -180
<< ndiff >>
rect -20 -195 30 -180
rect -20 -265 -5 -195
rect 15 -265 30 -195
rect -20 -280 30 -265
rect 45 -195 95 -180
rect 45 -265 60 -195
rect 80 -265 95 -195
rect 45 -280 95 -265
rect 110 -195 160 -180
rect 110 -265 125 -195
rect 145 -265 160 -195
rect 110 -280 160 -265
rect 230 -195 280 -180
rect 230 -265 245 -195
rect 265 -265 280 -195
rect 230 -280 280 -265
rect 295 -195 345 -180
rect 295 -265 310 -195
rect 330 -265 345 -195
rect 295 -280 345 -265
rect 360 -195 410 -180
rect 360 -265 375 -195
rect 395 -265 410 -195
rect 360 -280 410 -265
<< pdiff >>
rect -20 90 30 105
rect -20 20 -5 90
rect 15 20 30 90
rect -20 5 30 20
rect 65 90 115 105
rect 65 20 80 90
rect 100 20 115 90
rect 65 5 115 20
rect 150 90 200 105
rect 150 20 165 90
rect 185 20 200 90
rect 150 5 200 20
rect 230 90 280 105
rect 230 20 245 90
rect 265 20 280 90
rect 230 5 280 20
rect 315 90 365 105
rect 315 20 330 90
rect 350 20 365 90
rect 315 5 365 20
<< ndiffc >>
rect -5 -265 15 -195
rect 60 -265 80 -195
rect 125 -265 145 -195
rect 245 -265 265 -195
rect 310 -265 330 -195
rect 375 -265 395 -195
<< pdiffc >>
rect -5 20 15 90
rect 80 20 100 90
rect 165 20 185 90
rect 245 20 265 90
rect 330 20 350 90
<< psubdiff >>
rect -100 -195 -50 -180
rect -100 -265 -85 -195
rect -65 -265 -50 -195
rect -100 -280 -50 -265
<< nsubdiff >>
rect -100 90 -50 105
rect -100 20 -85 90
rect -65 20 -50 90
rect -100 5 -50 20
<< psubdiffcont >>
rect -85 -265 -65 -195
<< nsubdiffcont >>
rect -85 20 -65 90
<< poly >>
rect 110 150 150 160
rect 110 135 120 150
rect 30 130 120 135
rect 140 130 150 150
rect 30 120 150 130
rect 275 150 315 160
rect 275 130 285 150
rect 305 130 315 150
rect 275 120 315 130
rect 30 105 65 120
rect 115 105 150 120
rect 280 105 315 120
rect 30 -10 65 5
rect 115 -10 150 5
rect 280 -10 315 5
rect 30 -180 45 -165
rect 95 -180 110 -165
rect 280 -180 295 -165
rect 345 -180 360 -165
rect 30 -295 45 -280
rect 0 -305 45 -295
rect 0 -325 10 -305
rect 30 -325 45 -305
rect 0 -335 45 -325
rect 95 -295 110 -280
rect 280 -295 295 -280
rect 345 -295 360 -280
rect 95 -305 140 -295
rect 95 -325 110 -305
rect 130 -325 140 -305
rect 280 -305 360 -295
rect 280 -310 310 -305
rect 95 -335 140 -325
rect 300 -325 310 -310
rect 330 -310 360 -305
rect 330 -325 340 -310
rect 300 -335 340 -325
<< polycont >>
rect 120 130 140 150
rect 285 130 305 150
rect 10 -325 30 -305
rect 110 -325 130 -305
rect 310 -325 330 -305
<< locali >>
rect 110 150 150 160
rect 275 150 315 160
rect -5 130 120 150
rect 140 130 150 150
rect -5 100 15 130
rect 110 120 150 130
rect 170 130 285 150
rect 305 130 315 150
rect 170 100 190 130
rect 275 120 315 130
rect -95 90 -55 100
rect -95 20 -85 90
rect -65 20 -55 90
rect -95 10 -55 20
rect -15 90 25 100
rect -15 20 -5 90
rect 15 20 25 90
rect -15 10 25 20
rect 70 90 110 100
rect 70 20 80 90
rect 100 20 110 90
rect 70 10 110 20
rect 155 90 195 100
rect 155 20 165 90
rect 185 20 195 90
rect 155 10 195 20
rect 235 90 275 100
rect 235 20 245 90
rect 265 20 275 90
rect 235 10 275 20
rect 320 90 360 100
rect 320 20 330 90
rect 350 20 360 90
rect 320 10 360 20
rect -5 -185 15 10
rect 50 -105 90 -95
rect 50 -125 60 -105
rect 80 -125 90 -105
rect 165 -115 185 10
rect 330 -70 350 10
rect 330 -90 470 -70
rect 50 -135 90 -125
rect 125 -135 185 -115
rect 235 -105 275 -95
rect 235 -125 245 -105
rect 265 -125 275 -105
rect 235 -135 275 -125
rect 60 -185 80 -135
rect 125 -185 145 -135
rect 245 -185 265 -135
rect 375 -185 395 -90
rect -95 -195 -55 -185
rect -95 -265 -85 -195
rect -65 -265 -55 -195
rect -95 -275 -55 -265
rect -15 -195 25 -185
rect -15 -265 -5 -195
rect 15 -265 25 -195
rect -15 -275 25 -265
rect 50 -195 90 -185
rect 50 -265 60 -195
rect 80 -265 90 -195
rect 50 -275 90 -265
rect 115 -195 155 -185
rect 115 -265 125 -195
rect 145 -265 155 -195
rect 115 -275 155 -265
rect 235 -195 275 -185
rect 235 -265 245 -195
rect 265 -265 275 -195
rect 235 -275 275 -265
rect 300 -195 340 -185
rect 300 -265 310 -195
rect 330 -265 340 -195
rect 300 -275 340 -265
rect 365 -195 405 -185
rect 365 -265 375 -195
rect 395 -265 405 -195
rect 365 -275 405 -265
rect 0 -305 40 -295
rect 0 -325 10 -305
rect 30 -325 40 -305
rect 0 -335 40 -325
rect 100 -305 140 -295
rect 100 -325 110 -305
rect 130 -325 140 -305
rect 100 -335 140 -325
rect 300 -305 340 -295
rect 300 -325 310 -305
rect 330 -325 340 -305
rect 300 -335 340 -325
<< viali >>
rect -85 20 -65 90
rect 80 20 100 90
rect 245 20 265 90
rect 60 -125 80 -105
rect 245 -125 265 -105
rect -85 -265 -65 -195
rect 310 -265 330 -195
<< metal1 >>
rect -140 90 470 100
rect -140 20 -85 90
rect -65 20 80 90
rect 100 20 245 90
rect 265 20 470 90
rect -140 10 470 20
rect 50 -105 275 -95
rect 50 -125 60 -105
rect 80 -125 245 -105
rect 265 -125 275 -105
rect 50 -135 275 -125
rect -140 -195 470 -185
rect -140 -265 -85 -195
rect -65 -265 310 -195
rect 330 -265 470 -195
rect -140 -275 470 -265
<< labels >>
rlabel metal1 -140 55 -140 55 1 VP
port 1 n
rlabel metal1 -140 -235 -140 -235 7 VN
port 2 w
rlabel locali 20 -335 20 -335 5 Vin_Minus
port 3 s
rlabel locali 120 -335 120 -335 5 Vin_Plus
port 4 s
rlabel locali 320 -335 320 -335 5 V_Bias
port 5 s
rlabel locali 470 -80 470 -80 3 Vout
port 6 e
<< end >>
