magic
tech sky130A
timestamp 1657193500
<< nwell >>
rect -160 225 435 375
<< pmoslvt >>
rect 0 250 35 350
rect 165 250 200 350
rect 330 250 365 350
<< nmoslvt >>
rect 55 55 70 155
rect 120 55 135 155
rect 265 55 280 155
<< ndiff >>
rect 5 140 55 155
rect 5 70 20 140
rect 40 70 55 140
rect 5 55 55 70
rect 70 140 120 155
rect 70 70 85 140
rect 105 70 120 140
rect 70 55 120 70
rect 135 140 185 155
rect 135 70 150 140
rect 170 70 185 140
rect 135 55 185 70
rect 215 140 265 155
rect 215 70 230 140
rect 250 70 265 140
rect 215 55 265 70
rect 280 140 330 155
rect 280 70 295 140
rect 315 70 330 140
rect 280 55 330 70
<< pdiff >>
rect -50 335 0 350
rect -50 265 -35 335
rect -15 265 0 335
rect -50 250 0 265
rect 35 335 85 350
rect 35 265 50 335
rect 70 265 85 335
rect 35 250 85 265
rect 115 335 165 350
rect 115 265 130 335
rect 150 265 165 335
rect 115 250 165 265
rect 200 335 250 350
rect 200 265 215 335
rect 235 265 250 335
rect 200 250 250 265
rect 280 335 330 350
rect 280 265 295 335
rect 315 265 330 335
rect 280 250 330 265
rect 365 335 415 350
rect 365 265 380 335
rect 400 265 415 335
rect 365 250 415 265
<< ndiffc >>
rect 20 70 40 140
rect 85 70 105 140
rect 150 70 170 140
rect 230 70 250 140
rect 295 70 315 140
<< pdiffc >>
rect -35 265 -15 335
rect 50 265 70 335
rect 130 265 150 335
rect 215 265 235 335
rect 295 265 315 335
rect 380 265 400 335
<< psubdiff >>
rect -75 145 -25 155
rect -75 70 -60 145
rect -40 70 -25 145
rect -75 55 -25 70
<< nsubdiff >>
rect -130 340 -80 350
rect -130 265 -115 340
rect -95 265 -80 340
rect -130 250 -80 265
<< psubdiffcont >>
rect -60 70 -40 145
<< nsubdiffcont >>
rect -115 265 -95 340
<< poly >>
rect 0 350 35 365
rect 165 350 200 365
rect 330 350 365 365
rect 0 240 35 250
rect 165 240 200 250
rect 330 240 365 250
rect 0 225 70 240
rect 55 155 70 225
rect 120 225 200 240
rect 265 225 365 240
rect 120 155 135 225
rect 265 215 280 225
rect 240 205 280 215
rect 240 185 250 205
rect 270 185 280 205
rect 240 175 280 185
rect 265 155 280 175
rect 55 40 70 55
rect 120 40 135 55
rect 265 40 280 55
<< polycont >>
rect 250 185 270 205
<< locali >>
rect -125 340 -85 345
rect -125 265 -115 340
rect -95 265 -85 340
rect -125 255 -85 265
rect -45 335 -5 345
rect -45 265 -35 335
rect -15 265 -5 335
rect -45 255 -5 265
rect 40 335 80 345
rect 40 265 50 335
rect 70 265 80 335
rect 40 255 80 265
rect 120 335 160 345
rect 120 265 130 335
rect 150 265 160 335
rect 120 255 160 265
rect 205 335 245 345
rect 205 265 215 335
rect 235 265 245 335
rect 205 255 245 265
rect 285 335 325 345
rect 285 265 295 335
rect 315 265 325 335
rect 285 255 325 265
rect 370 335 410 345
rect 370 265 380 335
rect 400 265 410 335
rect 370 255 410 265
rect -35 205 -15 255
rect 130 205 150 255
rect 240 205 280 215
rect -35 185 250 205
rect 270 185 280 205
rect 20 150 40 185
rect 240 175 280 185
rect 300 205 320 255
rect 300 185 435 205
rect 300 150 320 185
rect -70 145 -30 150
rect -70 70 -60 145
rect -40 70 -30 145
rect -70 60 -30 70
rect 10 140 50 150
rect 10 70 20 140
rect 40 70 50 140
rect 10 60 50 70
rect 75 140 115 150
rect 75 70 85 140
rect 105 70 115 140
rect 75 60 115 70
rect 140 140 180 150
rect 140 70 150 140
rect 170 70 180 140
rect 140 60 180 70
rect 220 140 260 150
rect 220 70 230 140
rect 250 70 260 140
rect 220 60 260 70
rect 285 140 325 150
rect 285 70 295 140
rect 315 70 325 140
rect 285 60 325 70
<< viali >>
rect -115 265 -95 340
rect 50 265 70 335
rect 215 265 235 335
rect 380 265 400 335
rect -60 70 -40 145
rect 150 70 170 140
rect 230 70 250 140
<< metal1 >>
rect -160 340 435 345
rect -160 265 -115 340
rect -95 335 435 340
rect -95 265 50 335
rect 70 265 215 335
rect 235 265 380 335
rect 400 265 435 335
rect -160 255 435 265
rect -160 145 435 150
rect -160 70 -60 145
rect -40 140 435 145
rect -40 70 150 140
rect 170 70 230 140
rect 250 70 435 140
rect -160 60 435 70
<< end >>
