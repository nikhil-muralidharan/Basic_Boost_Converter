magic
tech sky130A
magscale 1 2
timestamp 1658393137
<< nwell >>
rect -250 -30 1290 240
<< pmoslvt >>
rect 60 10 130 200
rect 390 10 460 200
rect 730 10 800 200
rect 1070 10 1140 200
rect 1926 50 1996 240
rect 2256 50 2326 240
<< nmoslvt >>
rect 1956 -360 1986 -170
rect 2086 -360 2118 -170
rect 80 -620 110 -430
rect 390 -620 420 -430
rect 700 -620 730 -430
<< ndiff >>
rect -20 -460 80 -430
rect -20 -590 10 -460
rect 50 -590 80 -460
rect -20 -620 80 -590
rect 110 -460 210 -430
rect 110 -590 140 -460
rect 180 -590 210 -460
rect 110 -620 210 -590
rect 290 -460 390 -430
rect 290 -590 320 -460
rect 360 -590 390 -460
rect 290 -620 390 -590
rect 420 -460 520 -430
rect 420 -590 450 -460
rect 490 -590 520 -460
rect 420 -620 520 -590
rect 600 -460 700 -430
rect 600 -590 630 -460
rect 670 -590 700 -460
rect 600 -620 700 -590
rect 730 -460 830 -430
rect 730 -590 760 -460
rect 800 -590 830 -460
rect 730 -620 830 -590
<< pdiff >>
rect -40 170 60 200
rect -40 40 -10 170
rect 30 40 60 170
rect -40 10 60 40
rect 130 170 230 200
rect 130 40 160 170
rect 200 40 230 170
rect 130 10 230 40
rect 290 170 390 200
rect 290 40 320 170
rect 360 40 390 170
rect 290 10 390 40
rect 460 170 560 200
rect 460 40 490 170
rect 530 40 560 170
rect 460 10 560 40
rect 630 170 730 200
rect 630 40 660 170
rect 700 40 730 170
rect 630 10 730 40
rect 800 170 900 200
rect 800 40 830 170
rect 870 40 900 170
rect 800 10 900 40
rect 970 170 1070 200
rect 970 40 1000 170
rect 1040 40 1070 170
rect 970 10 1070 40
rect 1140 170 1240 200
rect 1140 40 1170 170
rect 1210 40 1240 170
rect 1140 10 1240 40
<< ndiffc >>
rect 10 -590 50 -460
rect 140 -590 180 -460
rect 320 -590 360 -460
rect 450 -590 490 -460
rect 630 -590 670 -460
rect 760 -590 800 -460
<< pdiffc >>
rect -10 40 30 170
rect 160 40 200 170
rect 320 40 360 170
rect 490 40 530 170
rect 660 40 700 170
rect 830 40 870 170
rect 1000 40 1040 170
rect 1170 40 1210 170
<< psubdiff >>
rect -200 -460 -100 -430
rect -200 -590 -170 -460
rect -130 -590 -100 -460
rect -200 -620 -100 -590
<< nsubdiff >>
rect -200 170 -100 200
rect -200 40 -170 170
rect -130 40 -100 170
rect -200 10 -100 40
<< psubdiffcont >>
rect -170 -590 -130 -460
<< nsubdiffcont >>
rect -170 40 -130 170
<< poly >>
rect 20 440 130 460
rect 20 400 40 440
rect 80 400 130 440
rect 20 380 130 400
rect 350 440 460 460
rect 350 400 370 440
rect 410 400 460 440
rect 350 380 460 400
rect 690 440 800 460
rect 690 400 710 440
rect 750 400 800 440
rect 690 380 800 400
rect 1030 440 1140 460
rect 1030 400 1050 440
rect 1090 400 1140 440
rect 1030 380 1140 400
rect 60 200 130 380
rect 390 200 460 380
rect 730 200 800 380
rect 1070 200 1140 380
rect 60 -30 130 10
rect 390 -30 460 10
rect 730 -30 800 10
rect 1070 -30 1140 10
rect -5 -270 75 -250
rect -5 -310 15 -270
rect 55 -290 75 -270
rect 55 -310 730 -290
rect -5 -320 730 -310
rect -5 -330 75 -320
rect 80 -410 420 -380
rect 80 -430 110 -410
rect 390 -430 420 -410
rect 700 -430 730 -320
rect 80 -725 110 -620
rect 390 -650 420 -620
rect 700 -650 730 -620
rect 80 -745 160 -725
rect 80 -785 100 -745
rect 140 -785 160 -745
rect 80 -805 160 -785
<< polycont >>
rect 40 400 80 440
rect 370 400 410 440
rect 710 400 750 440
rect 1050 400 1090 440
rect 15 -310 55 -270
rect 100 -785 140 -745
<< locali >>
rect 40 460 80 500
rect 370 460 410 500
rect 20 440 100 460
rect 20 400 40 440
rect 80 400 100 440
rect 20 380 100 400
rect 350 440 430 460
rect 350 400 370 440
rect 410 400 430 440
rect 350 380 430 400
rect 550 300 600 500
rect 710 460 750 500
rect 1050 460 1090 500
rect 690 440 770 460
rect 690 400 710 440
rect 750 400 770 440
rect 690 380 770 400
rect 1030 440 1110 460
rect 1030 400 1050 440
rect 1090 400 1110 440
rect 1030 380 1110 400
rect 160 260 1450 300
rect 160 190 200 260
rect 490 190 530 260
rect 830 190 880 260
rect 1170 190 1220 260
rect -190 170 -110 190
rect -190 40 -170 170
rect -130 40 -110 170
rect -190 20 -110 40
rect -30 170 50 190
rect -30 40 -10 170
rect 30 40 50 170
rect -30 20 50 40
rect 140 170 220 190
rect 140 40 160 170
rect 200 40 220 170
rect 140 20 220 40
rect 300 170 380 190
rect 300 40 320 170
rect 360 40 380 170
rect 300 20 380 40
rect 470 170 550 190
rect 470 40 490 170
rect 530 40 550 170
rect 470 20 550 40
rect 640 170 720 190
rect 640 40 660 170
rect 700 40 720 170
rect 640 20 720 40
rect 810 170 890 190
rect 810 40 830 170
rect 870 40 890 170
rect 810 20 890 40
rect 980 170 1060 190
rect 980 40 1000 170
rect 1040 40 1060 170
rect 980 20 1060 40
rect 1150 170 1230 190
rect 1150 40 1170 170
rect 1210 40 1230 170
rect 1150 20 1230 40
rect -10 -140 30 20
rect 320 -50 360 20
rect 660 -50 700 20
rect 320 -90 700 -50
rect 660 -130 700 -90
rect -10 -180 50 -140
rect 10 -250 50 -180
rect 610 -170 700 -130
rect 610 -220 650 -170
rect 1000 -210 1040 20
rect -5 -270 75 -250
rect -5 -310 15 -270
rect 55 -310 75 -270
rect -5 -330 75 -310
rect 140 -260 650 -220
rect 690 -250 1040 -210
rect 10 -440 50 -390
rect 140 -440 180 -260
rect 690 -300 730 -250
rect 450 -340 730 -300
rect 450 -440 490 -340
rect 1410 -360 1450 260
rect 760 -400 1540 -360
rect 760 -440 800 -400
rect 1500 -440 1660 -400
rect -190 -460 -110 -440
rect -190 -590 -170 -460
rect -130 -590 -110 -460
rect -190 -610 -110 -590
rect -10 -460 70 -440
rect -10 -590 10 -460
rect 50 -590 70 -460
rect -10 -610 70 -590
rect 120 -460 200 -440
rect 120 -590 140 -460
rect 180 -590 200 -460
rect 120 -610 200 -590
rect 300 -460 380 -440
rect 300 -590 320 -460
rect 360 -590 380 -460
rect 300 -610 380 -590
rect 430 -460 510 -440
rect 430 -590 450 -460
rect 490 -590 510 -460
rect 430 -610 510 -590
rect 610 -460 690 -440
rect 610 -590 630 -460
rect 670 -590 690 -460
rect 610 -610 690 -590
rect 740 -460 820 -440
rect 740 -590 760 -460
rect 800 -590 820 -460
rect 740 -610 820 -590
rect 10 -650 50 -610
rect -40 -690 50 -650
rect 140 -650 180 -610
rect 140 -690 260 -650
rect -40 -840 0 -690
rect 80 -740 160 -725
rect 220 -740 260 -690
rect 80 -745 260 -740
rect 80 -785 100 -745
rect 140 -780 260 -745
rect 140 -785 160 -780
rect 80 -805 160 -785
rect 320 -840 360 -610
rect 630 -840 670 -610
rect -40 -880 670 -840
<< viali >>
rect -170 40 -130 170
rect 160 40 200 170
rect 490 40 530 170
rect 830 40 870 170
rect 1170 40 1210 170
rect -170 -590 -130 -460
rect 10 -590 50 -460
rect 320 -590 360 -460
rect 630 -590 670 -460
<< metal1 >>
rect -250 170 1290 190
rect -250 40 -170 170
rect -130 40 160 170
rect 200 40 490 170
rect 530 40 830 170
rect 870 40 1170 170
rect 1210 40 1290 170
rect -250 20 1290 40
rect -250 -460 1290 -440
rect -250 -590 -170 -460
rect -130 -590 10 -460
rect 50 -590 320 -460
rect 360 -590 630 -460
rect 670 -590 1290 -460
rect -250 -610 1290 -590
use BUFFER  BUFFER_0
timestamp 1658392951
transform 1 0 2836 0 1 -200
box -1240 -260 -358 492
<< labels >>
rlabel space 2478 -90 2478 -90 3 Vout
port 4 e
rlabel locali 310 -880 310 -880 5 Gnd
port 6 s
rlabel locali 570 500 570 500 1 Idc
port 5 n
rlabel locali 60 500 60 500 1 Vref
port 7 n
rlabel locali 390 500 390 500 1 Vofb
port 8 n
rlabel locali 730 500 730 500 1 Vsen
port 9 n
rlabel locali 1070 500 1070 500 1 Vsen_DC
port 10 n
<< end >>
