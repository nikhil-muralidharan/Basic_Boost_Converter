magic
tech sky130A
timestamp 1657893085
<< nwell >>
rect -280 40 490 190
<< pmoslvt >>
rect -125 70 -90 170
rect 45 70 80 170
rect 215 70 250 170
rect 385 70 420 170
<< nmoslvt >>
rect -115 -85 -100 5
rect 45 -85 60 5
rect 205 -85 220 5
rect 365 -85 380 5
<< ndiff >>
rect -175 -5 -115 5
rect -175 -65 -155 -5
rect -135 -65 -115 -5
rect -175 -85 -115 -65
rect -100 -5 -45 5
rect -100 -65 -80 -5
rect -60 -65 -45 -5
rect -100 -85 -45 -65
rect -15 -5 45 5
rect -15 -65 5 -5
rect 25 -65 45 -5
rect -15 -85 45 -65
rect 60 -5 115 5
rect 60 -65 80 -5
rect 100 -65 115 -5
rect 60 -85 115 -65
rect 145 -5 205 5
rect 145 -65 165 -5
rect 185 -65 205 -5
rect 145 -85 205 -65
rect 220 -5 275 5
rect 220 -65 240 -5
rect 260 -65 275 -5
rect 220 -85 275 -65
rect 305 -5 365 5
rect 305 -65 325 -5
rect 345 -65 365 -5
rect 305 -85 365 -65
rect 380 -5 435 5
rect 380 -65 400 -5
rect 420 -65 435 -5
rect 380 -85 435 -65
<< pdiff >>
rect -180 155 -125 170
rect -180 85 -160 155
rect -140 85 -125 155
rect -180 70 -125 85
rect -90 155 -40 170
rect -90 85 -75 155
rect -55 85 -40 155
rect -90 70 -40 85
rect -10 155 45 170
rect -10 85 10 155
rect 30 85 45 155
rect -10 70 45 85
rect 80 155 130 170
rect 80 85 95 155
rect 115 85 130 155
rect 80 70 130 85
rect 160 155 215 170
rect 160 85 180 155
rect 200 85 215 155
rect 160 70 215 85
rect 250 155 300 170
rect 250 85 265 155
rect 285 85 300 155
rect 250 70 300 85
rect 330 155 385 170
rect 330 85 350 155
rect 370 85 385 155
rect 330 70 385 85
rect 420 155 470 170
rect 420 85 435 155
rect 455 85 470 155
rect 420 70 470 85
<< ndiffc >>
rect -155 -65 -135 -5
rect -80 -65 -60 -5
rect 5 -65 25 -5
rect 80 -65 100 -5
rect 165 -65 185 -5
rect 240 -65 260 -5
rect 325 -65 345 -5
rect 400 -65 420 -5
<< pdiffc >>
rect -160 85 -140 155
rect -75 85 -55 155
rect 10 85 30 155
rect 95 85 115 155
rect 180 85 200 155
rect 265 85 285 155
rect 350 85 370 155
rect 435 85 455 155
<< psubdiff >>
rect -255 -5 -205 5
rect -255 -65 -240 -5
rect -220 -65 -205 -5
rect -255 -85 -205 -65
<< nsubdiff >>
rect -260 155 -210 170
rect -260 85 -245 155
rect -225 85 -210 155
rect -260 70 -210 85
<< psubdiffcont >>
rect -240 -65 -220 -5
<< nsubdiffcont >>
rect -245 85 -225 155
<< poly >>
rect -125 170 -90 185
rect 45 170 80 185
rect 215 170 250 185
rect 385 170 420 185
rect -125 35 -90 70
rect -115 5 -100 35
rect 45 30 80 70
rect 215 35 250 70
rect 385 35 420 70
rect 45 5 60 30
rect 205 20 230 35
rect 365 30 420 35
rect 365 20 400 30
rect 205 5 220 20
rect 365 5 380 20
rect -115 -100 -100 -85
rect 45 -100 60 -85
rect 205 -100 220 -85
rect 365 -100 380 -85
rect -140 -110 -100 -100
rect -140 -130 -130 -110
rect -110 -130 -100 -110
rect -140 -140 -100 -130
rect 20 -110 60 -100
rect 20 -130 30 -110
rect 50 -130 60 -110
rect 20 -140 60 -130
rect 180 -110 220 -100
rect 180 -130 190 -110
rect 210 -130 220 -110
rect 180 -140 220 -130
rect 340 -110 380 -100
rect 340 -130 350 -110
rect 370 -130 380 -110
rect 340 -140 380 -130
<< polycont >>
rect -130 -130 -110 -110
rect 30 -130 50 -110
rect 190 -130 210 -110
rect 350 -130 370 -110
<< locali >>
rect -255 155 -215 165
rect -255 85 -245 155
rect -225 85 -215 155
rect -255 75 -215 85
rect -170 155 -130 165
rect -170 85 -160 155
rect -140 85 -130 155
rect -170 75 -130 85
rect -85 155 -45 165
rect -85 85 -75 155
rect -55 85 -45 155
rect -85 75 -45 85
rect 0 155 40 165
rect 0 85 10 155
rect 30 85 40 155
rect 0 75 40 85
rect 85 155 125 165
rect 85 85 95 155
rect 115 85 125 155
rect 85 75 125 85
rect 170 155 210 165
rect 170 85 180 155
rect 200 85 210 155
rect 170 75 210 85
rect 255 155 295 165
rect 255 85 265 155
rect 285 85 295 155
rect 255 75 295 85
rect 340 155 380 165
rect 340 85 350 155
rect 370 85 380 155
rect 340 75 380 85
rect 425 155 465 165
rect 425 85 435 155
rect 455 85 465 155
rect 425 75 465 85
rect -75 45 -50 75
rect 95 45 120 75
rect -75 25 120 45
rect 265 45 290 75
rect 435 45 460 75
rect 265 25 460 45
rect 85 0 105 25
rect 405 0 425 25
rect -250 -5 -210 0
rect -250 -65 -240 -5
rect -220 -65 -210 -5
rect -250 -75 -210 -65
rect -165 -5 -125 0
rect -165 -65 -155 -5
rect -135 -65 -125 -5
rect -165 -75 -125 -65
rect -90 -5 -50 0
rect -90 -65 -80 -5
rect -60 -65 -50 -5
rect -90 -75 -50 -65
rect -5 -5 35 0
rect -5 -65 5 -5
rect 25 -65 35 -5
rect -5 -75 35 -65
rect 70 -5 110 0
rect 70 -65 80 -5
rect 100 -65 110 -5
rect 70 -75 110 -65
rect 155 -5 195 0
rect 155 -65 165 -5
rect 185 -65 195 -5
rect 155 -75 195 -65
rect 230 -5 270 0
rect 230 -65 240 -5
rect 260 -65 270 -5
rect 230 -75 270 -65
rect 315 -5 355 0
rect 315 -65 325 -5
rect 345 -65 355 -5
rect 315 -75 355 -65
rect 390 -5 430 0
rect 390 -65 400 -5
rect 420 -65 430 -5
rect 390 -75 430 -65
rect -140 -110 -100 -100
rect -140 -130 -130 -110
rect -110 -130 -100 -110
rect -140 -140 -100 -130
rect 20 -110 60 -100
rect 20 -130 30 -110
rect 50 -130 60 -110
rect 20 -140 60 -130
rect 180 -110 220 -100
rect 180 -130 190 -110
rect 210 -130 220 -110
rect 180 -140 220 -130
rect 340 -110 380 -100
rect 340 -130 350 -110
rect 370 -130 380 -110
rect 340 -140 380 -130
<< viali >>
rect -245 85 -225 155
rect -160 85 -140 155
rect 10 85 30 155
rect 180 85 200 155
rect 350 85 370 155
rect -240 -65 -220 -5
rect -155 -65 -135 -5
rect 165 -65 185 -5
<< metal1 >>
rect -280 155 490 165
rect -280 85 -245 155
rect -225 85 -160 155
rect -140 85 10 155
rect 30 85 180 155
rect 200 85 350 155
rect 370 85 490 155
rect -280 75 490 85
rect -280 -5 490 0
rect -280 -65 -240 -5
rect -220 -65 -155 -5
rect -135 -65 165 -5
rect 185 -65 490 -5
rect -280 -75 490 -65
<< labels >>
rlabel metal1 -280 -40 -280 -40 7 GND
rlabel metal1 -280 110 -280 110 7 VDD
rlabel poly -110 25 -110 25 7 S
rlabel poly 215 20 215 20 7 R
rlabel poly 50 15 50 15 7 Q
rlabel poly 370 15 370 15 7 ZCD
<< end >>
