magic
tech sky130A
timestamp 1641706646
<< psubdiff >>
rect 8690 11475 8775 11490
rect 8690 11435 8705 11475
rect 8745 11435 8775 11475
rect 8690 11420 8775 11435
rect 10355 11475 10440 11490
rect 10355 11435 10385 11475
rect 10425 11435 10440 11475
rect 10355 11420 10440 11435
rect 13645 11475 13730 11490
rect 13645 11435 13660 11475
rect 13700 11435 13730 11475
rect 13645 11420 13730 11435
rect 15310 11475 15395 11490
rect 15310 11435 15340 11475
rect 15380 11435 15395 11475
rect 15310 11420 15395 11435
rect 18600 11475 18685 11490
rect 18600 11435 18615 11475
rect 18655 11435 18685 11475
rect 18600 11420 18685 11435
rect 20265 11475 20350 11490
rect 20265 11435 20295 11475
rect 20335 11435 20350 11475
rect 20265 11420 20350 11435
rect 23555 11475 23640 11490
rect 23555 11435 23570 11475
rect 23610 11435 23640 11475
rect 23555 11420 23640 11435
rect 25220 11475 25305 11490
rect 25220 11435 25250 11475
rect 25290 11435 25305 11475
rect 25220 11420 25305 11435
rect 28510 11475 28595 11490
rect 28510 11435 28525 11475
rect 28565 11435 28595 11475
rect 28510 11420 28595 11435
rect 30175 11475 30260 11490
rect 30175 11435 30205 11475
rect 30245 11435 30260 11475
rect 30175 11420 30260 11435
rect 33465 11475 33550 11490
rect 33465 11435 33480 11475
rect 33520 11435 33550 11475
rect 33465 11420 33550 11435
rect 35130 11475 35215 11490
rect 35130 11435 35160 11475
rect 35200 11435 35215 11475
rect 35130 11420 35215 11435
rect 38420 11475 38505 11490
rect 38420 11435 38435 11475
rect 38475 11435 38505 11475
rect 38420 11420 38505 11435
rect 40085 11475 40170 11490
rect 40085 11435 40115 11475
rect 40155 11435 40170 11475
rect 40085 11420 40170 11435
rect 43375 11475 43460 11490
rect 43375 11435 43390 11475
rect 43430 11435 43460 11475
rect 43375 11420 43460 11435
rect 45040 11475 45125 11490
rect 45040 11435 45070 11475
rect 45110 11435 45125 11475
rect 45040 11420 45125 11435
rect 48330 11475 48415 11490
rect 48330 11435 48345 11475
rect 48385 11435 48415 11475
rect 48330 11420 48415 11435
rect 49995 11475 50080 11490
rect 49995 11435 50025 11475
rect 50065 11435 50080 11475
rect 49995 11420 50080 11435
rect 53285 11475 53370 11490
rect 53285 11435 53300 11475
rect 53340 11435 53370 11475
rect 53285 11420 53370 11435
rect 54950 11475 55035 11490
rect 54950 11435 54980 11475
rect 55020 11435 55035 11475
rect 54950 11420 55035 11435
rect 58240 11475 58325 11490
rect 58240 11435 58255 11475
rect 58295 11435 58325 11475
rect 58240 11420 58325 11435
rect 59905 11475 59990 11490
rect 59905 11435 59935 11475
rect 59975 11435 59990 11475
rect 59905 11420 59990 11435
rect 63195 11475 63280 11490
rect 63195 11435 63210 11475
rect 63250 11435 63280 11475
rect 63195 11420 63280 11435
rect 64860 11475 64945 11490
rect 64860 11435 64890 11475
rect 64930 11435 64945 11475
rect 64860 11420 64945 11435
rect 68150 11475 68235 11490
rect 68150 11435 68165 11475
rect 68205 11435 68235 11475
rect 68150 11420 68235 11435
rect 69815 11475 69900 11490
rect 69815 11435 69845 11475
rect 69885 11435 69900 11475
rect 69815 11420 69900 11435
rect 73105 11475 73190 11490
rect 73105 11435 73120 11475
rect 73160 11435 73190 11475
rect 73105 11420 73190 11435
rect 74770 11475 74855 11490
rect 74770 11435 74800 11475
rect 74840 11435 74855 11475
rect 74770 11420 74855 11435
rect 8690 9555 8775 9570
rect 8690 9515 8705 9555
rect 8745 9515 8775 9555
rect 8690 9500 8775 9515
rect 10355 9555 10440 9570
rect 10355 9515 10385 9555
rect 10425 9515 10440 9555
rect 10355 9500 10440 9515
rect 13645 9555 13730 9570
rect 13645 9515 13660 9555
rect 13700 9515 13730 9555
rect 13645 9500 13730 9515
rect 15310 9555 15395 9570
rect 15310 9515 15340 9555
rect 15380 9515 15395 9555
rect 15310 9500 15395 9515
rect 18600 9555 18685 9570
rect 18600 9515 18615 9555
rect 18655 9515 18685 9555
rect 18600 9500 18685 9515
rect 20265 9555 20350 9570
rect 20265 9515 20295 9555
rect 20335 9515 20350 9555
rect 20265 9500 20350 9515
rect 23555 9555 23640 9570
rect 23555 9515 23570 9555
rect 23610 9515 23640 9555
rect 23555 9500 23640 9515
rect 25220 9555 25305 9570
rect 25220 9515 25250 9555
rect 25290 9515 25305 9555
rect 25220 9500 25305 9515
rect 28510 9555 28595 9570
rect 28510 9515 28525 9555
rect 28565 9515 28595 9555
rect 28510 9500 28595 9515
rect 30175 9555 30260 9570
rect 30175 9515 30205 9555
rect 30245 9515 30260 9555
rect 30175 9500 30260 9515
rect 33465 9555 33550 9570
rect 33465 9515 33480 9555
rect 33520 9515 33550 9555
rect 33465 9500 33550 9515
rect 35130 9555 35215 9570
rect 35130 9515 35160 9555
rect 35200 9515 35215 9555
rect 35130 9500 35215 9515
rect 38420 9555 38505 9570
rect 38420 9515 38435 9555
rect 38475 9515 38505 9555
rect 38420 9500 38505 9515
rect 40085 9555 40170 9570
rect 40085 9515 40115 9555
rect 40155 9515 40170 9555
rect 40085 9500 40170 9515
rect 43375 9555 43460 9570
rect 43375 9515 43390 9555
rect 43430 9515 43460 9555
rect 43375 9500 43460 9515
rect 45040 9555 45125 9570
rect 45040 9515 45070 9555
rect 45110 9515 45125 9555
rect 45040 9500 45125 9515
rect 48330 9555 48415 9570
rect 48330 9515 48345 9555
rect 48385 9515 48415 9555
rect 48330 9500 48415 9515
rect 49995 9555 50080 9570
rect 49995 9515 50025 9555
rect 50065 9515 50080 9555
rect 49995 9500 50080 9515
rect 53285 9555 53370 9570
rect 53285 9515 53300 9555
rect 53340 9515 53370 9555
rect 53285 9500 53370 9515
rect 54950 9555 55035 9570
rect 54950 9515 54980 9555
rect 55020 9515 55035 9555
rect 54950 9500 55035 9515
rect 58240 9555 58325 9570
rect 58240 9515 58255 9555
rect 58295 9515 58325 9555
rect 58240 9500 58325 9515
rect 59905 9555 59990 9570
rect 59905 9515 59935 9555
rect 59975 9515 59990 9555
rect 59905 9500 59990 9515
rect 63195 9555 63280 9570
rect 63195 9515 63210 9555
rect 63250 9515 63280 9555
rect 63195 9500 63280 9515
rect 64860 9555 64945 9570
rect 64860 9515 64890 9555
rect 64930 9515 64945 9555
rect 64860 9500 64945 9515
rect 68150 9555 68235 9570
rect 68150 9515 68165 9555
rect 68205 9515 68235 9555
rect 68150 9500 68235 9515
rect 69815 9555 69900 9570
rect 69815 9515 69845 9555
rect 69885 9515 69900 9555
rect 69815 9500 69900 9515
rect 73105 9555 73190 9570
rect 73105 9515 73120 9555
rect 73160 9515 73190 9555
rect 73105 9500 73190 9515
rect 74770 9555 74855 9570
rect 74770 9515 74800 9555
rect 74840 9515 74855 9555
rect 74770 9500 74855 9515
rect 5615 9270 5685 9285
rect 5615 9230 5630 9270
rect 5670 9230 5685 9270
rect 5615 9200 5685 9230
rect 6815 9270 6885 9285
rect 6815 9230 6830 9270
rect 6870 9230 6885 9270
rect 6815 9200 6885 9230
rect 7295 9270 7365 9285
rect 7295 9230 7310 9270
rect 7350 9230 7365 9270
rect 7295 9200 7365 9230
rect 8495 9270 8565 9285
rect 8495 9230 8510 9270
rect 8550 9230 8565 9270
rect 8495 9200 8565 9230
rect 10570 9270 10640 9285
rect 10570 9230 10585 9270
rect 10625 9230 10640 9270
rect 10570 9200 10640 9230
rect 11770 9270 11840 9285
rect 11770 9230 11785 9270
rect 11825 9230 11840 9270
rect 11770 9200 11840 9230
rect 12250 9270 12320 9285
rect 12250 9230 12265 9270
rect 12305 9230 12320 9270
rect 12250 9200 12320 9230
rect 13450 9270 13520 9285
rect 13450 9230 13465 9270
rect 13505 9230 13520 9270
rect 13450 9200 13520 9230
rect 15525 9270 15595 9285
rect 15525 9230 15540 9270
rect 15580 9230 15595 9270
rect 15525 9200 15595 9230
rect 16725 9270 16795 9285
rect 16725 9230 16740 9270
rect 16780 9230 16795 9270
rect 16725 9200 16795 9230
rect 17205 9270 17275 9285
rect 17205 9230 17220 9270
rect 17260 9230 17275 9270
rect 17205 9200 17275 9230
rect 18405 9270 18475 9285
rect 18405 9230 18420 9270
rect 18460 9230 18475 9270
rect 18405 9200 18475 9230
rect 20480 9270 20550 9285
rect 20480 9230 20495 9270
rect 20535 9230 20550 9270
rect 20480 9200 20550 9230
rect 21680 9270 21750 9285
rect 21680 9230 21695 9270
rect 21735 9230 21750 9270
rect 21680 9200 21750 9230
rect 22160 9270 22230 9285
rect 22160 9230 22175 9270
rect 22215 9230 22230 9270
rect 22160 9200 22230 9230
rect 23360 9270 23430 9285
rect 23360 9230 23375 9270
rect 23415 9230 23430 9270
rect 23360 9200 23430 9230
rect 25435 9270 25505 9285
rect 25435 9230 25450 9270
rect 25490 9230 25505 9270
rect 25435 9200 25505 9230
rect 26635 9270 26705 9285
rect 26635 9230 26650 9270
rect 26690 9230 26705 9270
rect 26635 9200 26705 9230
rect 27115 9270 27185 9285
rect 27115 9230 27130 9270
rect 27170 9230 27185 9270
rect 27115 9200 27185 9230
rect 28315 9270 28385 9285
rect 28315 9230 28330 9270
rect 28370 9230 28385 9270
rect 28315 9200 28385 9230
rect 30390 9270 30460 9285
rect 30390 9230 30405 9270
rect 30445 9230 30460 9270
rect 30390 9200 30460 9230
rect 31590 9270 31660 9285
rect 31590 9230 31605 9270
rect 31645 9230 31660 9270
rect 31590 9200 31660 9230
rect 32070 9270 32140 9285
rect 32070 9230 32085 9270
rect 32125 9230 32140 9270
rect 32070 9200 32140 9230
rect 33270 9270 33340 9285
rect 33270 9230 33285 9270
rect 33325 9230 33340 9270
rect 33270 9200 33340 9230
rect 35345 9270 35415 9285
rect 35345 9230 35360 9270
rect 35400 9230 35415 9270
rect 35345 9200 35415 9230
rect 36545 9270 36615 9285
rect 36545 9230 36560 9270
rect 36600 9230 36615 9270
rect 36545 9200 36615 9230
rect 37025 9270 37095 9285
rect 37025 9230 37040 9270
rect 37080 9230 37095 9270
rect 37025 9200 37095 9230
rect 38225 9270 38295 9285
rect 38225 9230 38240 9270
rect 38280 9230 38295 9270
rect 38225 9200 38295 9230
rect 40300 9270 40370 9285
rect 40300 9230 40315 9270
rect 40355 9230 40370 9270
rect 40300 9200 40370 9230
rect 41500 9270 41570 9285
rect 41500 9230 41515 9270
rect 41555 9230 41570 9270
rect 41500 9200 41570 9230
rect 41980 9270 42050 9285
rect 41980 9230 41995 9270
rect 42035 9230 42050 9270
rect 41980 9200 42050 9230
rect 43180 9270 43250 9285
rect 43180 9230 43195 9270
rect 43235 9230 43250 9270
rect 43180 9200 43250 9230
rect 45255 9270 45325 9285
rect 45255 9230 45270 9270
rect 45310 9230 45325 9270
rect 45255 9200 45325 9230
rect 46455 9270 46525 9285
rect 46455 9230 46470 9270
rect 46510 9230 46525 9270
rect 46455 9200 46525 9230
rect 46935 9270 47005 9285
rect 46935 9230 46950 9270
rect 46990 9230 47005 9270
rect 46935 9200 47005 9230
rect 48135 9270 48205 9285
rect 48135 9230 48150 9270
rect 48190 9230 48205 9270
rect 48135 9200 48205 9230
rect 50210 9270 50280 9285
rect 50210 9230 50225 9270
rect 50265 9230 50280 9270
rect 50210 9200 50280 9230
rect 51410 9270 51480 9285
rect 51410 9230 51425 9270
rect 51465 9230 51480 9270
rect 51410 9200 51480 9230
rect 51890 9270 51960 9285
rect 51890 9230 51905 9270
rect 51945 9230 51960 9270
rect 51890 9200 51960 9230
rect 53090 9270 53160 9285
rect 53090 9230 53105 9270
rect 53145 9230 53160 9270
rect 53090 9200 53160 9230
rect 55165 9270 55235 9285
rect 55165 9230 55180 9270
rect 55220 9230 55235 9270
rect 55165 9200 55235 9230
rect 56365 9270 56435 9285
rect 56365 9230 56380 9270
rect 56420 9230 56435 9270
rect 56365 9200 56435 9230
rect 56845 9270 56915 9285
rect 56845 9230 56860 9270
rect 56900 9230 56915 9270
rect 56845 9200 56915 9230
rect 58045 9270 58115 9285
rect 58045 9230 58060 9270
rect 58100 9230 58115 9270
rect 58045 9200 58115 9230
rect 60120 9270 60190 9285
rect 60120 9230 60135 9270
rect 60175 9230 60190 9270
rect 60120 9200 60190 9230
rect 61320 9270 61390 9285
rect 61320 9230 61335 9270
rect 61375 9230 61390 9270
rect 61320 9200 61390 9230
rect 61800 9270 61870 9285
rect 61800 9230 61815 9270
rect 61855 9230 61870 9270
rect 61800 9200 61870 9230
rect 63000 9270 63070 9285
rect 63000 9230 63015 9270
rect 63055 9230 63070 9270
rect 63000 9200 63070 9230
rect 65075 9270 65145 9285
rect 65075 9230 65090 9270
rect 65130 9230 65145 9270
rect 65075 9200 65145 9230
rect 66275 9270 66345 9285
rect 66275 9230 66290 9270
rect 66330 9230 66345 9270
rect 66275 9200 66345 9230
rect 66755 9270 66825 9285
rect 66755 9230 66770 9270
rect 66810 9230 66825 9270
rect 66755 9200 66825 9230
rect 67955 9270 68025 9285
rect 67955 9230 67970 9270
rect 68010 9230 68025 9270
rect 67955 9200 68025 9230
rect 70030 9270 70100 9285
rect 70030 9230 70045 9270
rect 70085 9230 70100 9270
rect 70030 9200 70100 9230
rect 71230 9270 71300 9285
rect 71230 9230 71245 9270
rect 71285 9230 71300 9270
rect 71230 9200 71300 9230
rect 71710 9270 71780 9285
rect 71710 9230 71725 9270
rect 71765 9230 71780 9270
rect 71710 9200 71780 9230
rect 72910 9270 72980 9285
rect 72910 9230 72925 9270
rect 72965 9230 72980 9270
rect 72910 9200 72980 9230
rect 74985 9270 75055 9285
rect 74985 9230 75000 9270
rect 75040 9230 75055 9270
rect 74985 9200 75055 9230
rect 76185 9270 76255 9285
rect 76185 9230 76200 9270
rect 76240 9230 76255 9270
rect 76185 9200 76255 9230
rect 76665 9270 76735 9285
rect 76665 9230 76680 9270
rect 76720 9230 76735 9270
rect 76665 9200 76735 9230
rect 77865 9270 77935 9285
rect 77865 9230 77880 9270
rect 77920 9230 77935 9270
rect 77865 9200 77935 9230
rect 5615 8640 5685 8670
rect 5615 8600 5630 8640
rect 5670 8600 5685 8640
rect 5615 8585 5685 8600
rect 6815 8640 6885 8670
rect 6815 8600 6830 8640
rect 6870 8600 6885 8640
rect 6815 8585 6885 8600
rect 7295 8640 7365 8670
rect 7295 8600 7310 8640
rect 7350 8600 7365 8640
rect 7295 8585 7365 8600
rect 8495 8640 8565 8670
rect 8495 8600 8510 8640
rect 8550 8600 8565 8640
rect 8495 8585 8565 8600
rect 10570 8640 10640 8670
rect 10570 8600 10585 8640
rect 10625 8600 10640 8640
rect 10570 8585 10640 8600
rect 11770 8640 11840 8670
rect 11770 8600 11785 8640
rect 11825 8600 11840 8640
rect 11770 8585 11840 8600
rect 12250 8640 12320 8670
rect 12250 8600 12265 8640
rect 12305 8600 12320 8640
rect 12250 8585 12320 8600
rect 13450 8640 13520 8670
rect 13450 8600 13465 8640
rect 13505 8600 13520 8640
rect 13450 8585 13520 8600
rect 15525 8640 15595 8670
rect 15525 8600 15540 8640
rect 15580 8600 15595 8640
rect 15525 8585 15595 8600
rect 16725 8640 16795 8670
rect 16725 8600 16740 8640
rect 16780 8600 16795 8640
rect 16725 8585 16795 8600
rect 17205 8640 17275 8670
rect 17205 8600 17220 8640
rect 17260 8600 17275 8640
rect 17205 8585 17275 8600
rect 18405 8640 18475 8670
rect 18405 8600 18420 8640
rect 18460 8600 18475 8640
rect 18405 8585 18475 8600
rect 20480 8640 20550 8670
rect 20480 8600 20495 8640
rect 20535 8600 20550 8640
rect 20480 8585 20550 8600
rect 21680 8640 21750 8670
rect 21680 8600 21695 8640
rect 21735 8600 21750 8640
rect 21680 8585 21750 8600
rect 22160 8640 22230 8670
rect 22160 8600 22175 8640
rect 22215 8600 22230 8640
rect 22160 8585 22230 8600
rect 23360 8640 23430 8670
rect 23360 8600 23375 8640
rect 23415 8600 23430 8640
rect 23360 8585 23430 8600
rect 25435 8640 25505 8670
rect 25435 8600 25450 8640
rect 25490 8600 25505 8640
rect 25435 8585 25505 8600
rect 26635 8640 26705 8670
rect 26635 8600 26650 8640
rect 26690 8600 26705 8640
rect 26635 8585 26705 8600
rect 27115 8640 27185 8670
rect 27115 8600 27130 8640
rect 27170 8600 27185 8640
rect 27115 8585 27185 8600
rect 28315 8640 28385 8670
rect 28315 8600 28330 8640
rect 28370 8600 28385 8640
rect 28315 8585 28385 8600
rect 30390 8640 30460 8670
rect 30390 8600 30405 8640
rect 30445 8600 30460 8640
rect 30390 8585 30460 8600
rect 31590 8640 31660 8670
rect 31590 8600 31605 8640
rect 31645 8600 31660 8640
rect 31590 8585 31660 8600
rect 32070 8640 32140 8670
rect 32070 8600 32085 8640
rect 32125 8600 32140 8640
rect 32070 8585 32140 8600
rect 33270 8640 33340 8670
rect 33270 8600 33285 8640
rect 33325 8600 33340 8640
rect 33270 8585 33340 8600
rect 35345 8640 35415 8670
rect 35345 8600 35360 8640
rect 35400 8600 35415 8640
rect 35345 8585 35415 8600
rect 36545 8640 36615 8670
rect 36545 8600 36560 8640
rect 36600 8600 36615 8640
rect 36545 8585 36615 8600
rect 37025 8640 37095 8670
rect 37025 8600 37040 8640
rect 37080 8600 37095 8640
rect 37025 8585 37095 8600
rect 38225 8640 38295 8670
rect 38225 8600 38240 8640
rect 38280 8600 38295 8640
rect 38225 8585 38295 8600
rect 40300 8640 40370 8670
rect 40300 8600 40315 8640
rect 40355 8600 40370 8640
rect 40300 8585 40370 8600
rect 41500 8640 41570 8670
rect 41500 8600 41515 8640
rect 41555 8600 41570 8640
rect 41500 8585 41570 8600
rect 41980 8640 42050 8670
rect 41980 8600 41995 8640
rect 42035 8600 42050 8640
rect 41980 8585 42050 8600
rect 43180 8640 43250 8670
rect 43180 8600 43195 8640
rect 43235 8600 43250 8640
rect 43180 8585 43250 8600
rect 45255 8640 45325 8670
rect 45255 8600 45270 8640
rect 45310 8600 45325 8640
rect 45255 8585 45325 8600
rect 46455 8640 46525 8670
rect 46455 8600 46470 8640
rect 46510 8600 46525 8640
rect 46455 8585 46525 8600
rect 46935 8640 47005 8670
rect 46935 8600 46950 8640
rect 46990 8600 47005 8640
rect 46935 8585 47005 8600
rect 48135 8640 48205 8670
rect 48135 8600 48150 8640
rect 48190 8600 48205 8640
rect 48135 8585 48205 8600
rect 50210 8640 50280 8670
rect 50210 8600 50225 8640
rect 50265 8600 50280 8640
rect 50210 8585 50280 8600
rect 51410 8640 51480 8670
rect 51410 8600 51425 8640
rect 51465 8600 51480 8640
rect 51410 8585 51480 8600
rect 51890 8640 51960 8670
rect 51890 8600 51905 8640
rect 51945 8600 51960 8640
rect 51890 8585 51960 8600
rect 53090 8640 53160 8670
rect 53090 8600 53105 8640
rect 53145 8600 53160 8640
rect 53090 8585 53160 8600
rect 55165 8640 55235 8670
rect 55165 8600 55180 8640
rect 55220 8600 55235 8640
rect 55165 8585 55235 8600
rect 56365 8640 56435 8670
rect 56365 8600 56380 8640
rect 56420 8600 56435 8640
rect 56365 8585 56435 8600
rect 56845 8640 56915 8670
rect 56845 8600 56860 8640
rect 56900 8600 56915 8640
rect 56845 8585 56915 8600
rect 58045 8640 58115 8670
rect 58045 8600 58060 8640
rect 58100 8600 58115 8640
rect 58045 8585 58115 8600
rect 60120 8640 60190 8670
rect 60120 8600 60135 8640
rect 60175 8600 60190 8640
rect 60120 8585 60190 8600
rect 61320 8640 61390 8670
rect 61320 8600 61335 8640
rect 61375 8600 61390 8640
rect 61320 8585 61390 8600
rect 61800 8640 61870 8670
rect 61800 8600 61815 8640
rect 61855 8600 61870 8640
rect 61800 8585 61870 8600
rect 63000 8640 63070 8670
rect 63000 8600 63015 8640
rect 63055 8600 63070 8640
rect 63000 8585 63070 8600
rect 65075 8640 65145 8670
rect 65075 8600 65090 8640
rect 65130 8600 65145 8640
rect 65075 8585 65145 8600
rect 66275 8640 66345 8670
rect 66275 8600 66290 8640
rect 66330 8600 66345 8640
rect 66275 8585 66345 8600
rect 66755 8640 66825 8670
rect 66755 8600 66770 8640
rect 66810 8600 66825 8640
rect 66755 8585 66825 8600
rect 67955 8640 68025 8670
rect 67955 8600 67970 8640
rect 68010 8600 68025 8640
rect 67955 8585 68025 8600
rect 70030 8640 70100 8670
rect 70030 8600 70045 8640
rect 70085 8600 70100 8640
rect 70030 8585 70100 8600
rect 71230 8640 71300 8670
rect 71230 8600 71245 8640
rect 71285 8600 71300 8640
rect 71230 8585 71300 8600
rect 71710 8640 71780 8670
rect 71710 8600 71725 8640
rect 71765 8600 71780 8640
rect 71710 8585 71780 8600
rect 72910 8640 72980 8670
rect 72910 8600 72925 8640
rect 72965 8600 72980 8640
rect 72910 8585 72980 8600
rect 74985 8640 75055 8670
rect 74985 8600 75000 8640
rect 75040 8600 75055 8640
rect 74985 8585 75055 8600
rect 76185 8640 76255 8670
rect 76185 8600 76200 8640
rect 76240 8600 76255 8640
rect 76185 8585 76255 8600
rect 76665 8640 76735 8670
rect 76665 8600 76680 8640
rect 76720 8600 76735 8640
rect 76665 8585 76735 8600
rect 77865 8640 77935 8670
rect 77865 8600 77880 8640
rect 77920 8600 77935 8640
rect 77865 8585 77935 8600
rect 8690 8400 8775 8415
rect 8690 8360 8705 8400
rect 8745 8360 8775 8400
rect 8690 8345 8775 8360
rect 10355 8400 10440 8415
rect 10355 8360 10385 8400
rect 10425 8360 10440 8400
rect 10355 8345 10440 8360
rect 13645 8400 13730 8415
rect 13645 8360 13660 8400
rect 13700 8360 13730 8400
rect 13645 8345 13730 8360
rect 15310 8400 15395 8415
rect 15310 8360 15340 8400
rect 15380 8360 15395 8400
rect 15310 8345 15395 8360
rect 18600 8400 18685 8415
rect 18600 8360 18615 8400
rect 18655 8360 18685 8400
rect 18600 8345 18685 8360
rect 20265 8400 20350 8415
rect 20265 8360 20295 8400
rect 20335 8360 20350 8400
rect 20265 8345 20350 8360
rect 23555 8400 23640 8415
rect 23555 8360 23570 8400
rect 23610 8360 23640 8400
rect 23555 8345 23640 8360
rect 25220 8400 25305 8415
rect 25220 8360 25250 8400
rect 25290 8360 25305 8400
rect 25220 8345 25305 8360
rect 28510 8400 28595 8415
rect 28510 8360 28525 8400
rect 28565 8360 28595 8400
rect 28510 8345 28595 8360
rect 30175 8400 30260 8415
rect 30175 8360 30205 8400
rect 30245 8360 30260 8400
rect 30175 8345 30260 8360
rect 33465 8400 33550 8415
rect 33465 8360 33480 8400
rect 33520 8360 33550 8400
rect 33465 8345 33550 8360
rect 35130 8400 35215 8415
rect 35130 8360 35160 8400
rect 35200 8360 35215 8400
rect 35130 8345 35215 8360
rect 38420 8400 38505 8415
rect 38420 8360 38435 8400
rect 38475 8360 38505 8400
rect 38420 8345 38505 8360
rect 40085 8400 40170 8415
rect 40085 8360 40115 8400
rect 40155 8360 40170 8400
rect 40085 8345 40170 8360
rect 43375 8400 43460 8415
rect 43375 8360 43390 8400
rect 43430 8360 43460 8400
rect 43375 8345 43460 8360
rect 45040 8400 45125 8415
rect 45040 8360 45070 8400
rect 45110 8360 45125 8400
rect 45040 8345 45125 8360
rect 48330 8400 48415 8415
rect 48330 8360 48345 8400
rect 48385 8360 48415 8400
rect 48330 8345 48415 8360
rect 49995 8400 50080 8415
rect 49995 8360 50025 8400
rect 50065 8360 50080 8400
rect 49995 8345 50080 8360
rect 53285 8400 53370 8415
rect 53285 8360 53300 8400
rect 53340 8360 53370 8400
rect 53285 8345 53370 8360
rect 54950 8400 55035 8415
rect 54950 8360 54980 8400
rect 55020 8360 55035 8400
rect 54950 8345 55035 8360
rect 58240 8400 58325 8415
rect 58240 8360 58255 8400
rect 58295 8360 58325 8400
rect 58240 8345 58325 8360
rect 59905 8400 59990 8415
rect 59905 8360 59935 8400
rect 59975 8360 59990 8400
rect 59905 8345 59990 8360
rect 63195 8400 63280 8415
rect 63195 8360 63210 8400
rect 63250 8360 63280 8400
rect 63195 8345 63280 8360
rect 64860 8400 64945 8415
rect 64860 8360 64890 8400
rect 64930 8360 64945 8400
rect 64860 8345 64945 8360
rect 68150 8400 68235 8415
rect 68150 8360 68165 8400
rect 68205 8360 68235 8400
rect 68150 8345 68235 8360
rect 69815 8400 69900 8415
rect 69815 8360 69845 8400
rect 69885 8360 69900 8400
rect 69815 8345 69900 8360
rect 73105 8400 73190 8415
rect 73105 8360 73120 8400
rect 73160 8360 73190 8400
rect 73105 8345 73190 8360
rect 74770 8400 74855 8415
rect 74770 8360 74800 8400
rect 74840 8360 74855 8400
rect 74770 8345 74855 8360
rect 8690 6480 8775 6495
rect 8690 6440 8705 6480
rect 8745 6440 8775 6480
rect 8690 6425 8775 6440
rect 10355 6480 10440 6495
rect 10355 6440 10385 6480
rect 10425 6440 10440 6480
rect 10355 6425 10440 6440
rect 13645 6480 13730 6495
rect 13645 6440 13660 6480
rect 13700 6440 13730 6480
rect 13645 6425 13730 6440
rect 15310 6480 15395 6495
rect 15310 6440 15340 6480
rect 15380 6440 15395 6480
rect 15310 6425 15395 6440
rect 18600 6480 18685 6495
rect 18600 6440 18615 6480
rect 18655 6440 18685 6480
rect 18600 6425 18685 6440
rect 20265 6480 20350 6495
rect 20265 6440 20295 6480
rect 20335 6440 20350 6480
rect 20265 6425 20350 6440
rect 23555 6480 23640 6495
rect 23555 6440 23570 6480
rect 23610 6440 23640 6480
rect 23555 6425 23640 6440
rect 25220 6480 25305 6495
rect 25220 6440 25250 6480
rect 25290 6440 25305 6480
rect 25220 6425 25305 6440
rect 28510 6480 28595 6495
rect 28510 6440 28525 6480
rect 28565 6440 28595 6480
rect 28510 6425 28595 6440
rect 30175 6480 30260 6495
rect 30175 6440 30205 6480
rect 30245 6440 30260 6480
rect 30175 6425 30260 6440
rect 33465 6480 33550 6495
rect 33465 6440 33480 6480
rect 33520 6440 33550 6480
rect 33465 6425 33550 6440
rect 35130 6480 35215 6495
rect 35130 6440 35160 6480
rect 35200 6440 35215 6480
rect 35130 6425 35215 6440
rect 38420 6480 38505 6495
rect 38420 6440 38435 6480
rect 38475 6440 38505 6480
rect 38420 6425 38505 6440
rect 40085 6480 40170 6495
rect 40085 6440 40115 6480
rect 40155 6440 40170 6480
rect 40085 6425 40170 6440
rect 43375 6480 43460 6495
rect 43375 6440 43390 6480
rect 43430 6440 43460 6480
rect 43375 6425 43460 6440
rect 45040 6480 45125 6495
rect 45040 6440 45070 6480
rect 45110 6440 45125 6480
rect 45040 6425 45125 6440
rect 48330 6480 48415 6495
rect 48330 6440 48345 6480
rect 48385 6440 48415 6480
rect 48330 6425 48415 6440
rect 49995 6480 50080 6495
rect 49995 6440 50025 6480
rect 50065 6440 50080 6480
rect 49995 6425 50080 6440
rect 53285 6480 53370 6495
rect 53285 6440 53300 6480
rect 53340 6440 53370 6480
rect 53285 6425 53370 6440
rect 54950 6480 55035 6495
rect 54950 6440 54980 6480
rect 55020 6440 55035 6480
rect 54950 6425 55035 6440
rect 58240 6480 58325 6495
rect 58240 6440 58255 6480
rect 58295 6440 58325 6480
rect 58240 6425 58325 6440
rect 59905 6480 59990 6495
rect 59905 6440 59935 6480
rect 59975 6440 59990 6480
rect 59905 6425 59990 6440
rect 63195 6480 63280 6495
rect 63195 6440 63210 6480
rect 63250 6440 63280 6480
rect 63195 6425 63280 6440
rect 64860 6480 64945 6495
rect 64860 6440 64890 6480
rect 64930 6440 64945 6480
rect 64860 6425 64945 6440
rect 68150 6480 68235 6495
rect 68150 6440 68165 6480
rect 68205 6440 68235 6480
rect 68150 6425 68235 6440
rect 69815 6480 69900 6495
rect 69815 6440 69845 6480
rect 69885 6440 69900 6480
rect 69815 6425 69900 6440
rect 73105 6480 73190 6495
rect 73105 6440 73120 6480
rect 73160 6440 73190 6480
rect 73105 6425 73190 6440
rect 74770 6480 74855 6495
rect 74770 6440 74800 6480
rect 74840 6440 74855 6480
rect 74770 6425 74855 6440
rect 5615 6195 5685 6210
rect 5615 6155 5630 6195
rect 5670 6155 5685 6195
rect 5615 6125 5685 6155
rect 6815 6195 6885 6210
rect 6815 6155 6830 6195
rect 6870 6155 6885 6195
rect 6815 6125 6885 6155
rect 7295 6195 7365 6210
rect 7295 6155 7310 6195
rect 7350 6155 7365 6195
rect 7295 6125 7365 6155
rect 8495 6195 8565 6210
rect 8495 6155 8510 6195
rect 8550 6155 8565 6195
rect 8495 6125 8565 6155
rect 10570 6195 10640 6210
rect 10570 6155 10585 6195
rect 10625 6155 10640 6195
rect 10570 6125 10640 6155
rect 11770 6195 11840 6210
rect 11770 6155 11785 6195
rect 11825 6155 11840 6195
rect 11770 6125 11840 6155
rect 12250 6195 12320 6210
rect 12250 6155 12265 6195
rect 12305 6155 12320 6195
rect 12250 6125 12320 6155
rect 13450 6195 13520 6210
rect 13450 6155 13465 6195
rect 13505 6155 13520 6195
rect 13450 6125 13520 6155
rect 15525 6195 15595 6210
rect 15525 6155 15540 6195
rect 15580 6155 15595 6195
rect 15525 6125 15595 6155
rect 16725 6195 16795 6210
rect 16725 6155 16740 6195
rect 16780 6155 16795 6195
rect 16725 6125 16795 6155
rect 17205 6195 17275 6210
rect 17205 6155 17220 6195
rect 17260 6155 17275 6195
rect 17205 6125 17275 6155
rect 18405 6195 18475 6210
rect 18405 6155 18420 6195
rect 18460 6155 18475 6195
rect 18405 6125 18475 6155
rect 20480 6195 20550 6210
rect 20480 6155 20495 6195
rect 20535 6155 20550 6195
rect 20480 6125 20550 6155
rect 21680 6195 21750 6210
rect 21680 6155 21695 6195
rect 21735 6155 21750 6195
rect 21680 6125 21750 6155
rect 22160 6195 22230 6210
rect 22160 6155 22175 6195
rect 22215 6155 22230 6195
rect 22160 6125 22230 6155
rect 23360 6195 23430 6210
rect 23360 6155 23375 6195
rect 23415 6155 23430 6195
rect 23360 6125 23430 6155
rect 25435 6195 25505 6210
rect 25435 6155 25450 6195
rect 25490 6155 25505 6195
rect 25435 6125 25505 6155
rect 26635 6195 26705 6210
rect 26635 6155 26650 6195
rect 26690 6155 26705 6195
rect 26635 6125 26705 6155
rect 27115 6195 27185 6210
rect 27115 6155 27130 6195
rect 27170 6155 27185 6195
rect 27115 6125 27185 6155
rect 28315 6195 28385 6210
rect 28315 6155 28330 6195
rect 28370 6155 28385 6195
rect 28315 6125 28385 6155
rect 30390 6195 30460 6210
rect 30390 6155 30405 6195
rect 30445 6155 30460 6195
rect 30390 6125 30460 6155
rect 31590 6195 31660 6210
rect 31590 6155 31605 6195
rect 31645 6155 31660 6195
rect 31590 6125 31660 6155
rect 32070 6195 32140 6210
rect 32070 6155 32085 6195
rect 32125 6155 32140 6195
rect 32070 6125 32140 6155
rect 33270 6195 33340 6210
rect 33270 6155 33285 6195
rect 33325 6155 33340 6195
rect 33270 6125 33340 6155
rect 35345 6195 35415 6210
rect 35345 6155 35360 6195
rect 35400 6155 35415 6195
rect 35345 6125 35415 6155
rect 36545 6195 36615 6210
rect 36545 6155 36560 6195
rect 36600 6155 36615 6195
rect 36545 6125 36615 6155
rect 37025 6195 37095 6210
rect 37025 6155 37040 6195
rect 37080 6155 37095 6195
rect 37025 6125 37095 6155
rect 38225 6195 38295 6210
rect 38225 6155 38240 6195
rect 38280 6155 38295 6195
rect 38225 6125 38295 6155
rect 40300 6195 40370 6210
rect 40300 6155 40315 6195
rect 40355 6155 40370 6195
rect 40300 6125 40370 6155
rect 41500 6195 41570 6210
rect 41500 6155 41515 6195
rect 41555 6155 41570 6195
rect 41500 6125 41570 6155
rect 41980 6195 42050 6210
rect 41980 6155 41995 6195
rect 42035 6155 42050 6195
rect 41980 6125 42050 6155
rect 43180 6195 43250 6210
rect 43180 6155 43195 6195
rect 43235 6155 43250 6195
rect 43180 6125 43250 6155
rect 45255 6195 45325 6210
rect 45255 6155 45270 6195
rect 45310 6155 45325 6195
rect 45255 6125 45325 6155
rect 46455 6195 46525 6210
rect 46455 6155 46470 6195
rect 46510 6155 46525 6195
rect 46455 6125 46525 6155
rect 46935 6195 47005 6210
rect 46935 6155 46950 6195
rect 46990 6155 47005 6195
rect 46935 6125 47005 6155
rect 48135 6195 48205 6210
rect 48135 6155 48150 6195
rect 48190 6155 48205 6195
rect 48135 6125 48205 6155
rect 50210 6195 50280 6210
rect 50210 6155 50225 6195
rect 50265 6155 50280 6195
rect 50210 6125 50280 6155
rect 51410 6195 51480 6210
rect 51410 6155 51425 6195
rect 51465 6155 51480 6195
rect 51410 6125 51480 6155
rect 51890 6195 51960 6210
rect 51890 6155 51905 6195
rect 51945 6155 51960 6195
rect 51890 6125 51960 6155
rect 53090 6195 53160 6210
rect 53090 6155 53105 6195
rect 53145 6155 53160 6195
rect 53090 6125 53160 6155
rect 55165 6195 55235 6210
rect 55165 6155 55180 6195
rect 55220 6155 55235 6195
rect 55165 6125 55235 6155
rect 56365 6195 56435 6210
rect 56365 6155 56380 6195
rect 56420 6155 56435 6195
rect 56365 6125 56435 6155
rect 56845 6195 56915 6210
rect 56845 6155 56860 6195
rect 56900 6155 56915 6195
rect 56845 6125 56915 6155
rect 58045 6195 58115 6210
rect 58045 6155 58060 6195
rect 58100 6155 58115 6195
rect 58045 6125 58115 6155
rect 60120 6195 60190 6210
rect 60120 6155 60135 6195
rect 60175 6155 60190 6195
rect 60120 6125 60190 6155
rect 61320 6195 61390 6210
rect 61320 6155 61335 6195
rect 61375 6155 61390 6195
rect 61320 6125 61390 6155
rect 61800 6195 61870 6210
rect 61800 6155 61815 6195
rect 61855 6155 61870 6195
rect 61800 6125 61870 6155
rect 63000 6195 63070 6210
rect 63000 6155 63015 6195
rect 63055 6155 63070 6195
rect 63000 6125 63070 6155
rect 65075 6195 65145 6210
rect 65075 6155 65090 6195
rect 65130 6155 65145 6195
rect 65075 6125 65145 6155
rect 66275 6195 66345 6210
rect 66275 6155 66290 6195
rect 66330 6155 66345 6195
rect 66275 6125 66345 6155
rect 66755 6195 66825 6210
rect 66755 6155 66770 6195
rect 66810 6155 66825 6195
rect 66755 6125 66825 6155
rect 67955 6195 68025 6210
rect 67955 6155 67970 6195
rect 68010 6155 68025 6195
rect 67955 6125 68025 6155
rect 70030 6195 70100 6210
rect 70030 6155 70045 6195
rect 70085 6155 70100 6195
rect 70030 6125 70100 6155
rect 71230 6195 71300 6210
rect 71230 6155 71245 6195
rect 71285 6155 71300 6195
rect 71230 6125 71300 6155
rect 71710 6195 71780 6210
rect 71710 6155 71725 6195
rect 71765 6155 71780 6195
rect 71710 6125 71780 6155
rect 72910 6195 72980 6210
rect 72910 6155 72925 6195
rect 72965 6155 72980 6195
rect 72910 6125 72980 6155
rect 74985 6195 75055 6210
rect 74985 6155 75000 6195
rect 75040 6155 75055 6195
rect 74985 6125 75055 6155
rect 76185 6195 76255 6210
rect 76185 6155 76200 6195
rect 76240 6155 76255 6195
rect 76185 6125 76255 6155
rect 76665 6195 76735 6210
rect 76665 6155 76680 6195
rect 76720 6155 76735 6195
rect 76665 6125 76735 6155
rect 77865 6195 77935 6210
rect 77865 6155 77880 6195
rect 77920 6155 77935 6195
rect 77865 6125 77935 6155
rect 5615 5565 5685 5595
rect 5615 5525 5630 5565
rect 5670 5525 5685 5565
rect 5615 5510 5685 5525
rect 6815 5565 6885 5595
rect 6815 5525 6830 5565
rect 6870 5525 6885 5565
rect 6815 5510 6885 5525
rect 7295 5565 7365 5595
rect 7295 5525 7310 5565
rect 7350 5525 7365 5565
rect 7295 5510 7365 5525
rect 8495 5565 8565 5595
rect 8495 5525 8510 5565
rect 8550 5525 8565 5565
rect 8495 5510 8565 5525
rect 10570 5565 10640 5595
rect 10570 5525 10585 5565
rect 10625 5525 10640 5565
rect 10570 5510 10640 5525
rect 11770 5565 11840 5595
rect 11770 5525 11785 5565
rect 11825 5525 11840 5565
rect 11770 5510 11840 5525
rect 12250 5565 12320 5595
rect 12250 5525 12265 5565
rect 12305 5525 12320 5565
rect 12250 5510 12320 5525
rect 13450 5565 13520 5595
rect 13450 5525 13465 5565
rect 13505 5525 13520 5565
rect 13450 5510 13520 5525
rect 15525 5565 15595 5595
rect 15525 5525 15540 5565
rect 15580 5525 15595 5565
rect 15525 5510 15595 5525
rect 16725 5565 16795 5595
rect 16725 5525 16740 5565
rect 16780 5525 16795 5565
rect 16725 5510 16795 5525
rect 17205 5565 17275 5595
rect 17205 5525 17220 5565
rect 17260 5525 17275 5565
rect 17205 5510 17275 5525
rect 18405 5565 18475 5595
rect 18405 5525 18420 5565
rect 18460 5525 18475 5565
rect 18405 5510 18475 5525
rect 20480 5565 20550 5595
rect 20480 5525 20495 5565
rect 20535 5525 20550 5565
rect 20480 5510 20550 5525
rect 21680 5565 21750 5595
rect 21680 5525 21695 5565
rect 21735 5525 21750 5565
rect 21680 5510 21750 5525
rect 22160 5565 22230 5595
rect 22160 5525 22175 5565
rect 22215 5525 22230 5565
rect 22160 5510 22230 5525
rect 23360 5565 23430 5595
rect 23360 5525 23375 5565
rect 23415 5525 23430 5565
rect 23360 5510 23430 5525
rect 25435 5565 25505 5595
rect 25435 5525 25450 5565
rect 25490 5525 25505 5565
rect 25435 5510 25505 5525
rect 26635 5565 26705 5595
rect 26635 5525 26650 5565
rect 26690 5525 26705 5565
rect 26635 5510 26705 5525
rect 27115 5565 27185 5595
rect 27115 5525 27130 5565
rect 27170 5525 27185 5565
rect 27115 5510 27185 5525
rect 28315 5565 28385 5595
rect 28315 5525 28330 5565
rect 28370 5525 28385 5565
rect 28315 5510 28385 5525
rect 30390 5565 30460 5595
rect 30390 5525 30405 5565
rect 30445 5525 30460 5565
rect 30390 5510 30460 5525
rect 31590 5565 31660 5595
rect 31590 5525 31605 5565
rect 31645 5525 31660 5565
rect 31590 5510 31660 5525
rect 32070 5565 32140 5595
rect 32070 5525 32085 5565
rect 32125 5525 32140 5565
rect 32070 5510 32140 5525
rect 33270 5565 33340 5595
rect 33270 5525 33285 5565
rect 33325 5525 33340 5565
rect 33270 5510 33340 5525
rect 35345 5565 35415 5595
rect 35345 5525 35360 5565
rect 35400 5525 35415 5565
rect 35345 5510 35415 5525
rect 36545 5565 36615 5595
rect 36545 5525 36560 5565
rect 36600 5525 36615 5565
rect 36545 5510 36615 5525
rect 37025 5565 37095 5595
rect 37025 5525 37040 5565
rect 37080 5525 37095 5565
rect 37025 5510 37095 5525
rect 38225 5565 38295 5595
rect 38225 5525 38240 5565
rect 38280 5525 38295 5565
rect 38225 5510 38295 5525
rect 40300 5565 40370 5595
rect 40300 5525 40315 5565
rect 40355 5525 40370 5565
rect 40300 5510 40370 5525
rect 41500 5565 41570 5595
rect 41500 5525 41515 5565
rect 41555 5525 41570 5565
rect 41500 5510 41570 5525
rect 41980 5565 42050 5595
rect 41980 5525 41995 5565
rect 42035 5525 42050 5565
rect 41980 5510 42050 5525
rect 43180 5565 43250 5595
rect 43180 5525 43195 5565
rect 43235 5525 43250 5565
rect 43180 5510 43250 5525
rect 45255 5565 45325 5595
rect 45255 5525 45270 5565
rect 45310 5525 45325 5565
rect 45255 5510 45325 5525
rect 46455 5565 46525 5595
rect 46455 5525 46470 5565
rect 46510 5525 46525 5565
rect 46455 5510 46525 5525
rect 46935 5565 47005 5595
rect 46935 5525 46950 5565
rect 46990 5525 47005 5565
rect 46935 5510 47005 5525
rect 48135 5565 48205 5595
rect 48135 5525 48150 5565
rect 48190 5525 48205 5565
rect 48135 5510 48205 5525
rect 50210 5565 50280 5595
rect 50210 5525 50225 5565
rect 50265 5525 50280 5565
rect 50210 5510 50280 5525
rect 51410 5565 51480 5595
rect 51410 5525 51425 5565
rect 51465 5525 51480 5565
rect 51410 5510 51480 5525
rect 51890 5565 51960 5595
rect 51890 5525 51905 5565
rect 51945 5525 51960 5565
rect 51890 5510 51960 5525
rect 53090 5565 53160 5595
rect 53090 5525 53105 5565
rect 53145 5525 53160 5565
rect 53090 5510 53160 5525
rect 55165 5565 55235 5595
rect 55165 5525 55180 5565
rect 55220 5525 55235 5565
rect 55165 5510 55235 5525
rect 56365 5565 56435 5595
rect 56365 5525 56380 5565
rect 56420 5525 56435 5565
rect 56365 5510 56435 5525
rect 56845 5565 56915 5595
rect 56845 5525 56860 5565
rect 56900 5525 56915 5565
rect 56845 5510 56915 5525
rect 58045 5565 58115 5595
rect 58045 5525 58060 5565
rect 58100 5525 58115 5565
rect 58045 5510 58115 5525
rect 60120 5565 60190 5595
rect 60120 5525 60135 5565
rect 60175 5525 60190 5565
rect 60120 5510 60190 5525
rect 61320 5565 61390 5595
rect 61320 5525 61335 5565
rect 61375 5525 61390 5565
rect 61320 5510 61390 5525
rect 61800 5565 61870 5595
rect 61800 5525 61815 5565
rect 61855 5525 61870 5565
rect 61800 5510 61870 5525
rect 63000 5565 63070 5595
rect 63000 5525 63015 5565
rect 63055 5525 63070 5565
rect 63000 5510 63070 5525
rect 65075 5565 65145 5595
rect 65075 5525 65090 5565
rect 65130 5525 65145 5565
rect 65075 5510 65145 5525
rect 66275 5565 66345 5595
rect 66275 5525 66290 5565
rect 66330 5525 66345 5565
rect 66275 5510 66345 5525
rect 66755 5565 66825 5595
rect 66755 5525 66770 5565
rect 66810 5525 66825 5565
rect 66755 5510 66825 5525
rect 67955 5565 68025 5595
rect 67955 5525 67970 5565
rect 68010 5525 68025 5565
rect 67955 5510 68025 5525
rect 70030 5565 70100 5595
rect 70030 5525 70045 5565
rect 70085 5525 70100 5565
rect 70030 5510 70100 5525
rect 71230 5565 71300 5595
rect 71230 5525 71245 5565
rect 71285 5525 71300 5565
rect 71230 5510 71300 5525
rect 71710 5565 71780 5595
rect 71710 5525 71725 5565
rect 71765 5525 71780 5565
rect 71710 5510 71780 5525
rect 72910 5565 72980 5595
rect 72910 5525 72925 5565
rect 72965 5525 72980 5565
rect 72910 5510 72980 5525
rect 74985 5565 75055 5595
rect 74985 5525 75000 5565
rect 75040 5525 75055 5565
rect 74985 5510 75055 5525
rect 76185 5565 76255 5595
rect 76185 5525 76200 5565
rect 76240 5525 76255 5565
rect 76185 5510 76255 5525
rect 76665 5565 76735 5595
rect 76665 5525 76680 5565
rect 76720 5525 76735 5565
rect 76665 5510 76735 5525
rect 77865 5565 77935 5595
rect 77865 5525 77880 5565
rect 77920 5525 77935 5565
rect 77865 5510 77935 5525
rect 8690 5325 8775 5340
rect 8690 5285 8705 5325
rect 8745 5285 8775 5325
rect 8690 5270 8775 5285
rect 10355 5325 10440 5340
rect 10355 5285 10385 5325
rect 10425 5285 10440 5325
rect 10355 5270 10440 5285
rect 13645 5325 13730 5340
rect 13645 5285 13660 5325
rect 13700 5285 13730 5325
rect 13645 5270 13730 5285
rect 15310 5325 15395 5340
rect 15310 5285 15340 5325
rect 15380 5285 15395 5325
rect 15310 5270 15395 5285
rect 18600 5325 18685 5340
rect 18600 5285 18615 5325
rect 18655 5285 18685 5325
rect 18600 5270 18685 5285
rect 20265 5325 20350 5340
rect 20265 5285 20295 5325
rect 20335 5285 20350 5325
rect 20265 5270 20350 5285
rect 23555 5325 23640 5340
rect 23555 5285 23570 5325
rect 23610 5285 23640 5325
rect 23555 5270 23640 5285
rect 25220 5325 25305 5340
rect 25220 5285 25250 5325
rect 25290 5285 25305 5325
rect 25220 5270 25305 5285
rect 28510 5325 28595 5340
rect 28510 5285 28525 5325
rect 28565 5285 28595 5325
rect 28510 5270 28595 5285
rect 30175 5325 30260 5340
rect 30175 5285 30205 5325
rect 30245 5285 30260 5325
rect 30175 5270 30260 5285
rect 33465 5325 33550 5340
rect 33465 5285 33480 5325
rect 33520 5285 33550 5325
rect 33465 5270 33550 5285
rect 35130 5325 35215 5340
rect 35130 5285 35160 5325
rect 35200 5285 35215 5325
rect 35130 5270 35215 5285
rect 38420 5325 38505 5340
rect 38420 5285 38435 5325
rect 38475 5285 38505 5325
rect 38420 5270 38505 5285
rect 40085 5325 40170 5340
rect 40085 5285 40115 5325
rect 40155 5285 40170 5325
rect 40085 5270 40170 5285
rect 43375 5325 43460 5340
rect 43375 5285 43390 5325
rect 43430 5285 43460 5325
rect 43375 5270 43460 5285
rect 45040 5325 45125 5340
rect 45040 5285 45070 5325
rect 45110 5285 45125 5325
rect 45040 5270 45125 5285
rect 48330 5325 48415 5340
rect 48330 5285 48345 5325
rect 48385 5285 48415 5325
rect 48330 5270 48415 5285
rect 49995 5325 50080 5340
rect 49995 5285 50025 5325
rect 50065 5285 50080 5325
rect 49995 5270 50080 5285
rect 53285 5325 53370 5340
rect 53285 5285 53300 5325
rect 53340 5285 53370 5325
rect 53285 5270 53370 5285
rect 54950 5325 55035 5340
rect 54950 5285 54980 5325
rect 55020 5285 55035 5325
rect 54950 5270 55035 5285
rect 58240 5325 58325 5340
rect 58240 5285 58255 5325
rect 58295 5285 58325 5325
rect 58240 5270 58325 5285
rect 59905 5325 59990 5340
rect 59905 5285 59935 5325
rect 59975 5285 59990 5325
rect 59905 5270 59990 5285
rect 63195 5325 63280 5340
rect 63195 5285 63210 5325
rect 63250 5285 63280 5325
rect 63195 5270 63280 5285
rect 64860 5325 64945 5340
rect 64860 5285 64890 5325
rect 64930 5285 64945 5325
rect 64860 5270 64945 5285
rect 68150 5325 68235 5340
rect 68150 5285 68165 5325
rect 68205 5285 68235 5325
rect 68150 5270 68235 5285
rect 69815 5325 69900 5340
rect 69815 5285 69845 5325
rect 69885 5285 69900 5325
rect 69815 5270 69900 5285
rect 73105 5325 73190 5340
rect 73105 5285 73120 5325
rect 73160 5285 73190 5325
rect 73105 5270 73190 5285
rect 74770 5325 74855 5340
rect 74770 5285 74800 5325
rect 74840 5285 74855 5325
rect 74770 5270 74855 5285
rect 8690 3405 8775 3420
rect 8690 3365 8705 3405
rect 8745 3365 8775 3405
rect 8690 3350 8775 3365
rect 10355 3405 10440 3420
rect 10355 3365 10385 3405
rect 10425 3365 10440 3405
rect 10355 3350 10440 3365
rect 13645 3405 13730 3420
rect 13645 3365 13660 3405
rect 13700 3365 13730 3405
rect 13645 3350 13730 3365
rect 15310 3405 15395 3420
rect 15310 3365 15340 3405
rect 15380 3365 15395 3405
rect 15310 3350 15395 3365
rect 18600 3405 18685 3420
rect 18600 3365 18615 3405
rect 18655 3365 18685 3405
rect 18600 3350 18685 3365
rect 20265 3405 20350 3420
rect 20265 3365 20295 3405
rect 20335 3365 20350 3405
rect 20265 3350 20350 3365
rect 23555 3405 23640 3420
rect 23555 3365 23570 3405
rect 23610 3365 23640 3405
rect 23555 3350 23640 3365
rect 25220 3405 25305 3420
rect 25220 3365 25250 3405
rect 25290 3365 25305 3405
rect 25220 3350 25305 3365
rect 28510 3405 28595 3420
rect 28510 3365 28525 3405
rect 28565 3365 28595 3405
rect 28510 3350 28595 3365
rect 30175 3405 30260 3420
rect 30175 3365 30205 3405
rect 30245 3365 30260 3405
rect 30175 3350 30260 3365
rect 33465 3405 33550 3420
rect 33465 3365 33480 3405
rect 33520 3365 33550 3405
rect 33465 3350 33550 3365
rect 35130 3405 35215 3420
rect 35130 3365 35160 3405
rect 35200 3365 35215 3405
rect 35130 3350 35215 3365
rect 38420 3405 38505 3420
rect 38420 3365 38435 3405
rect 38475 3365 38505 3405
rect 38420 3350 38505 3365
rect 40085 3405 40170 3420
rect 40085 3365 40115 3405
rect 40155 3365 40170 3405
rect 40085 3350 40170 3365
rect 43375 3405 43460 3420
rect 43375 3365 43390 3405
rect 43430 3365 43460 3405
rect 43375 3350 43460 3365
rect 45040 3405 45125 3420
rect 45040 3365 45070 3405
rect 45110 3365 45125 3405
rect 45040 3350 45125 3365
rect 48330 3405 48415 3420
rect 48330 3365 48345 3405
rect 48385 3365 48415 3405
rect 48330 3350 48415 3365
rect 49995 3405 50080 3420
rect 49995 3365 50025 3405
rect 50065 3365 50080 3405
rect 49995 3350 50080 3365
rect 53285 3405 53370 3420
rect 53285 3365 53300 3405
rect 53340 3365 53370 3405
rect 53285 3350 53370 3365
rect 54950 3405 55035 3420
rect 54950 3365 54980 3405
rect 55020 3365 55035 3405
rect 54950 3350 55035 3365
rect 58240 3405 58325 3420
rect 58240 3365 58255 3405
rect 58295 3365 58325 3405
rect 58240 3350 58325 3365
rect 59905 3405 59990 3420
rect 59905 3365 59935 3405
rect 59975 3365 59990 3405
rect 59905 3350 59990 3365
rect 63195 3405 63280 3420
rect 63195 3365 63210 3405
rect 63250 3365 63280 3405
rect 63195 3350 63280 3365
rect 64860 3405 64945 3420
rect 64860 3365 64890 3405
rect 64930 3365 64945 3405
rect 64860 3350 64945 3365
rect 68150 3405 68235 3420
rect 68150 3365 68165 3405
rect 68205 3365 68235 3405
rect 68150 3350 68235 3365
rect 69815 3405 69900 3420
rect 69815 3365 69845 3405
rect 69885 3365 69900 3405
rect 69815 3350 69900 3365
rect 73105 3405 73190 3420
rect 73105 3365 73120 3405
rect 73160 3365 73190 3405
rect 73105 3350 73190 3365
rect 74770 3405 74855 3420
rect 74770 3365 74800 3405
rect 74840 3365 74855 3405
rect 74770 3350 74855 3365
rect 660 3120 730 3135
rect 660 3080 675 3120
rect 715 3080 730 3120
rect 660 3050 730 3080
rect 5615 3120 5685 3135
rect 5615 3080 5630 3120
rect 5670 3080 5685 3120
rect 5615 3050 5685 3080
rect 6815 3120 6885 3135
rect 6815 3080 6830 3120
rect 6870 3080 6885 3120
rect 6815 3050 6885 3080
rect 7295 3120 7365 3135
rect 7295 3080 7310 3120
rect 7350 3080 7365 3120
rect 7295 3050 7365 3080
rect 8495 3120 8565 3135
rect 8495 3080 8510 3120
rect 8550 3080 8565 3120
rect 8495 3050 8565 3080
rect 10570 3120 10640 3135
rect 10570 3080 10585 3120
rect 10625 3080 10640 3120
rect 10570 3050 10640 3080
rect 11770 3120 11840 3135
rect 11770 3080 11785 3120
rect 11825 3080 11840 3120
rect 11770 3050 11840 3080
rect 12250 3120 12320 3135
rect 12250 3080 12265 3120
rect 12305 3080 12320 3120
rect 12250 3050 12320 3080
rect 13450 3120 13520 3135
rect 13450 3080 13465 3120
rect 13505 3080 13520 3120
rect 13450 3050 13520 3080
rect 15525 3120 15595 3135
rect 15525 3080 15540 3120
rect 15580 3080 15595 3120
rect 15525 3050 15595 3080
rect 16725 3120 16795 3135
rect 16725 3080 16740 3120
rect 16780 3080 16795 3120
rect 16725 3050 16795 3080
rect 17205 3120 17275 3135
rect 17205 3080 17220 3120
rect 17260 3080 17275 3120
rect 17205 3050 17275 3080
rect 18405 3120 18475 3135
rect 18405 3080 18420 3120
rect 18460 3080 18475 3120
rect 18405 3050 18475 3080
rect 20480 3120 20550 3135
rect 20480 3080 20495 3120
rect 20535 3080 20550 3120
rect 20480 3050 20550 3080
rect 21680 3120 21750 3135
rect 21680 3080 21695 3120
rect 21735 3080 21750 3120
rect 21680 3050 21750 3080
rect 22160 3120 22230 3135
rect 22160 3080 22175 3120
rect 22215 3080 22230 3120
rect 22160 3050 22230 3080
rect 23360 3120 23430 3135
rect 23360 3080 23375 3120
rect 23415 3080 23430 3120
rect 23360 3050 23430 3080
rect 25435 3120 25505 3135
rect 25435 3080 25450 3120
rect 25490 3080 25505 3120
rect 25435 3050 25505 3080
rect 26635 3120 26705 3135
rect 26635 3080 26650 3120
rect 26690 3080 26705 3120
rect 26635 3050 26705 3080
rect 27115 3120 27185 3135
rect 27115 3080 27130 3120
rect 27170 3080 27185 3120
rect 27115 3050 27185 3080
rect 28315 3120 28385 3135
rect 28315 3080 28330 3120
rect 28370 3080 28385 3120
rect 28315 3050 28385 3080
rect 30390 3120 30460 3135
rect 30390 3080 30405 3120
rect 30445 3080 30460 3120
rect 30390 3050 30460 3080
rect 31590 3120 31660 3135
rect 31590 3080 31605 3120
rect 31645 3080 31660 3120
rect 31590 3050 31660 3080
rect 32070 3120 32140 3135
rect 32070 3080 32085 3120
rect 32125 3080 32140 3120
rect 32070 3050 32140 3080
rect 33270 3120 33340 3135
rect 33270 3080 33285 3120
rect 33325 3080 33340 3120
rect 33270 3050 33340 3080
rect 35345 3120 35415 3135
rect 35345 3080 35360 3120
rect 35400 3080 35415 3120
rect 35345 3050 35415 3080
rect 36545 3120 36615 3135
rect 36545 3080 36560 3120
rect 36600 3080 36615 3120
rect 36545 3050 36615 3080
rect 37025 3120 37095 3135
rect 37025 3080 37040 3120
rect 37080 3080 37095 3120
rect 37025 3050 37095 3080
rect 38225 3120 38295 3135
rect 38225 3080 38240 3120
rect 38280 3080 38295 3120
rect 38225 3050 38295 3080
rect 40300 3120 40370 3135
rect 40300 3080 40315 3120
rect 40355 3080 40370 3120
rect 40300 3050 40370 3080
rect 41500 3120 41570 3135
rect 41500 3080 41515 3120
rect 41555 3080 41570 3120
rect 41500 3050 41570 3080
rect 41980 3120 42050 3135
rect 41980 3080 41995 3120
rect 42035 3080 42050 3120
rect 41980 3050 42050 3080
rect 43180 3120 43250 3135
rect 43180 3080 43195 3120
rect 43235 3080 43250 3120
rect 43180 3050 43250 3080
rect 45255 3120 45325 3135
rect 45255 3080 45270 3120
rect 45310 3080 45325 3120
rect 45255 3050 45325 3080
rect 46455 3120 46525 3135
rect 46455 3080 46470 3120
rect 46510 3080 46525 3120
rect 46455 3050 46525 3080
rect 46935 3120 47005 3135
rect 46935 3080 46950 3120
rect 46990 3080 47005 3120
rect 46935 3050 47005 3080
rect 48135 3120 48205 3135
rect 48135 3080 48150 3120
rect 48190 3080 48205 3120
rect 48135 3050 48205 3080
rect 50210 3120 50280 3135
rect 50210 3080 50225 3120
rect 50265 3080 50280 3120
rect 50210 3050 50280 3080
rect 51410 3120 51480 3135
rect 51410 3080 51425 3120
rect 51465 3080 51480 3120
rect 51410 3050 51480 3080
rect 51890 3120 51960 3135
rect 51890 3080 51905 3120
rect 51945 3080 51960 3120
rect 51890 3050 51960 3080
rect 53090 3120 53160 3135
rect 53090 3080 53105 3120
rect 53145 3080 53160 3120
rect 53090 3050 53160 3080
rect 55165 3120 55235 3135
rect 55165 3080 55180 3120
rect 55220 3080 55235 3120
rect 55165 3050 55235 3080
rect 56365 3120 56435 3135
rect 56365 3080 56380 3120
rect 56420 3080 56435 3120
rect 56365 3050 56435 3080
rect 56845 3120 56915 3135
rect 56845 3080 56860 3120
rect 56900 3080 56915 3120
rect 56845 3050 56915 3080
rect 58045 3120 58115 3135
rect 58045 3080 58060 3120
rect 58100 3080 58115 3120
rect 58045 3050 58115 3080
rect 60120 3120 60190 3135
rect 60120 3080 60135 3120
rect 60175 3080 60190 3120
rect 60120 3050 60190 3080
rect 61320 3120 61390 3135
rect 61320 3080 61335 3120
rect 61375 3080 61390 3120
rect 61320 3050 61390 3080
rect 61800 3120 61870 3135
rect 61800 3080 61815 3120
rect 61855 3080 61870 3120
rect 61800 3050 61870 3080
rect 63000 3120 63070 3135
rect 63000 3080 63015 3120
rect 63055 3080 63070 3120
rect 63000 3050 63070 3080
rect 65075 3120 65145 3135
rect 65075 3080 65090 3120
rect 65130 3080 65145 3120
rect 65075 3050 65145 3080
rect 66275 3120 66345 3135
rect 66275 3080 66290 3120
rect 66330 3080 66345 3120
rect 66275 3050 66345 3080
rect 66755 3120 66825 3135
rect 66755 3080 66770 3120
rect 66810 3080 66825 3120
rect 66755 3050 66825 3080
rect 67955 3120 68025 3135
rect 67955 3080 67970 3120
rect 68010 3080 68025 3120
rect 67955 3050 68025 3080
rect 70030 3120 70100 3135
rect 70030 3080 70045 3120
rect 70085 3080 70100 3120
rect 70030 3050 70100 3080
rect 71230 3120 71300 3135
rect 71230 3080 71245 3120
rect 71285 3080 71300 3120
rect 71230 3050 71300 3080
rect 71710 3120 71780 3135
rect 71710 3080 71725 3120
rect 71765 3080 71780 3120
rect 71710 3050 71780 3080
rect 72910 3120 72980 3135
rect 72910 3080 72925 3120
rect 72965 3080 72980 3120
rect 72910 3050 72980 3080
rect 74985 3120 75055 3135
rect 74985 3080 75000 3120
rect 75040 3080 75055 3120
rect 74985 3050 75055 3080
rect 76185 3120 76255 3135
rect 76185 3080 76200 3120
rect 76240 3080 76255 3120
rect 76185 3050 76255 3080
rect 76665 3120 76735 3135
rect 76665 3080 76680 3120
rect 76720 3080 76735 3120
rect 76665 3050 76735 3080
rect 77865 3120 77935 3135
rect 77865 3080 77880 3120
rect 77920 3080 77935 3120
rect 77865 3050 77935 3080
rect 660 2490 730 2520
rect 660 2450 675 2490
rect 715 2450 730 2490
rect 660 2435 730 2450
rect 5615 2490 5685 2520
rect 5615 2450 5630 2490
rect 5670 2450 5685 2490
rect 5615 2435 5685 2450
rect 6815 2490 6885 2520
rect 6815 2450 6830 2490
rect 6870 2450 6885 2490
rect 6815 2435 6885 2450
rect 7295 2490 7365 2520
rect 7295 2450 7310 2490
rect 7350 2450 7365 2490
rect 7295 2435 7365 2450
rect 8495 2490 8565 2520
rect 8495 2450 8510 2490
rect 8550 2450 8565 2490
rect 8495 2435 8565 2450
rect 10570 2490 10640 2520
rect 10570 2450 10585 2490
rect 10625 2450 10640 2490
rect 10570 2435 10640 2450
rect 11770 2490 11840 2520
rect 11770 2450 11785 2490
rect 11825 2450 11840 2490
rect 11770 2435 11840 2450
rect 12250 2490 12320 2520
rect 12250 2450 12265 2490
rect 12305 2450 12320 2490
rect 12250 2435 12320 2450
rect 13450 2490 13520 2520
rect 13450 2450 13465 2490
rect 13505 2450 13520 2490
rect 13450 2435 13520 2450
rect 15525 2490 15595 2520
rect 15525 2450 15540 2490
rect 15580 2450 15595 2490
rect 15525 2435 15595 2450
rect 16725 2490 16795 2520
rect 16725 2450 16740 2490
rect 16780 2450 16795 2490
rect 16725 2435 16795 2450
rect 17205 2490 17275 2520
rect 17205 2450 17220 2490
rect 17260 2450 17275 2490
rect 17205 2435 17275 2450
rect 18405 2490 18475 2520
rect 18405 2450 18420 2490
rect 18460 2450 18475 2490
rect 18405 2435 18475 2450
rect 20480 2490 20550 2520
rect 20480 2450 20495 2490
rect 20535 2450 20550 2490
rect 20480 2435 20550 2450
rect 21680 2490 21750 2520
rect 21680 2450 21695 2490
rect 21735 2450 21750 2490
rect 21680 2435 21750 2450
rect 22160 2490 22230 2520
rect 22160 2450 22175 2490
rect 22215 2450 22230 2490
rect 22160 2435 22230 2450
rect 23360 2490 23430 2520
rect 23360 2450 23375 2490
rect 23415 2450 23430 2490
rect 23360 2435 23430 2450
rect 25435 2490 25505 2520
rect 25435 2450 25450 2490
rect 25490 2450 25505 2490
rect 25435 2435 25505 2450
rect 26635 2490 26705 2520
rect 26635 2450 26650 2490
rect 26690 2450 26705 2490
rect 26635 2435 26705 2450
rect 27115 2490 27185 2520
rect 27115 2450 27130 2490
rect 27170 2450 27185 2490
rect 27115 2435 27185 2450
rect 28315 2490 28385 2520
rect 28315 2450 28330 2490
rect 28370 2450 28385 2490
rect 28315 2435 28385 2450
rect 30390 2490 30460 2520
rect 30390 2450 30405 2490
rect 30445 2450 30460 2490
rect 30390 2435 30460 2450
rect 31590 2490 31660 2520
rect 31590 2450 31605 2490
rect 31645 2450 31660 2490
rect 31590 2435 31660 2450
rect 32070 2490 32140 2520
rect 32070 2450 32085 2490
rect 32125 2450 32140 2490
rect 32070 2435 32140 2450
rect 33270 2490 33340 2520
rect 33270 2450 33285 2490
rect 33325 2450 33340 2490
rect 33270 2435 33340 2450
rect 35345 2490 35415 2520
rect 35345 2450 35360 2490
rect 35400 2450 35415 2490
rect 35345 2435 35415 2450
rect 36545 2490 36615 2520
rect 36545 2450 36560 2490
rect 36600 2450 36615 2490
rect 36545 2435 36615 2450
rect 37025 2490 37095 2520
rect 37025 2450 37040 2490
rect 37080 2450 37095 2490
rect 37025 2435 37095 2450
rect 38225 2490 38295 2520
rect 38225 2450 38240 2490
rect 38280 2450 38295 2490
rect 38225 2435 38295 2450
rect 40300 2490 40370 2520
rect 40300 2450 40315 2490
rect 40355 2450 40370 2490
rect 40300 2435 40370 2450
rect 41500 2490 41570 2520
rect 41500 2450 41515 2490
rect 41555 2450 41570 2490
rect 41500 2435 41570 2450
rect 41980 2490 42050 2520
rect 41980 2450 41995 2490
rect 42035 2450 42050 2490
rect 41980 2435 42050 2450
rect 43180 2490 43250 2520
rect 43180 2450 43195 2490
rect 43235 2450 43250 2490
rect 43180 2435 43250 2450
rect 45255 2490 45325 2520
rect 45255 2450 45270 2490
rect 45310 2450 45325 2490
rect 45255 2435 45325 2450
rect 46455 2490 46525 2520
rect 46455 2450 46470 2490
rect 46510 2450 46525 2490
rect 46455 2435 46525 2450
rect 46935 2490 47005 2520
rect 46935 2450 46950 2490
rect 46990 2450 47005 2490
rect 46935 2435 47005 2450
rect 48135 2490 48205 2520
rect 48135 2450 48150 2490
rect 48190 2450 48205 2490
rect 48135 2435 48205 2450
rect 50210 2490 50280 2520
rect 50210 2450 50225 2490
rect 50265 2450 50280 2490
rect 50210 2435 50280 2450
rect 51410 2490 51480 2520
rect 51410 2450 51425 2490
rect 51465 2450 51480 2490
rect 51410 2435 51480 2450
rect 51890 2490 51960 2520
rect 51890 2450 51905 2490
rect 51945 2450 51960 2490
rect 51890 2435 51960 2450
rect 53090 2490 53160 2520
rect 53090 2450 53105 2490
rect 53145 2450 53160 2490
rect 53090 2435 53160 2450
rect 55165 2490 55235 2520
rect 55165 2450 55180 2490
rect 55220 2450 55235 2490
rect 55165 2435 55235 2450
rect 56365 2490 56435 2520
rect 56365 2450 56380 2490
rect 56420 2450 56435 2490
rect 56365 2435 56435 2450
rect 56845 2490 56915 2520
rect 56845 2450 56860 2490
rect 56900 2450 56915 2490
rect 56845 2435 56915 2450
rect 58045 2490 58115 2520
rect 58045 2450 58060 2490
rect 58100 2450 58115 2490
rect 58045 2435 58115 2450
rect 60120 2490 60190 2520
rect 60120 2450 60135 2490
rect 60175 2450 60190 2490
rect 60120 2435 60190 2450
rect 61320 2490 61390 2520
rect 61320 2450 61335 2490
rect 61375 2450 61390 2490
rect 61320 2435 61390 2450
rect 61800 2490 61870 2520
rect 61800 2450 61815 2490
rect 61855 2450 61870 2490
rect 61800 2435 61870 2450
rect 63000 2490 63070 2520
rect 63000 2450 63015 2490
rect 63055 2450 63070 2490
rect 63000 2435 63070 2450
rect 65075 2490 65145 2520
rect 65075 2450 65090 2490
rect 65130 2450 65145 2490
rect 65075 2435 65145 2450
rect 66275 2490 66345 2520
rect 66275 2450 66290 2490
rect 66330 2450 66345 2490
rect 66275 2435 66345 2450
rect 66755 2490 66825 2520
rect 66755 2450 66770 2490
rect 66810 2450 66825 2490
rect 66755 2435 66825 2450
rect 67955 2490 68025 2520
rect 67955 2450 67970 2490
rect 68010 2450 68025 2490
rect 67955 2435 68025 2450
rect 70030 2490 70100 2520
rect 70030 2450 70045 2490
rect 70085 2450 70100 2490
rect 70030 2435 70100 2450
rect 71230 2490 71300 2520
rect 71230 2450 71245 2490
rect 71285 2450 71300 2490
rect 71230 2435 71300 2450
rect 71710 2490 71780 2520
rect 71710 2450 71725 2490
rect 71765 2450 71780 2490
rect 71710 2435 71780 2450
rect 72910 2490 72980 2520
rect 72910 2450 72925 2490
rect 72965 2450 72980 2490
rect 72910 2435 72980 2450
rect 74985 2490 75055 2520
rect 74985 2450 75000 2490
rect 75040 2450 75055 2490
rect 74985 2435 75055 2450
rect 76185 2490 76255 2520
rect 76185 2450 76200 2490
rect 76240 2450 76255 2490
rect 76185 2435 76255 2450
rect 76665 2490 76735 2520
rect 76665 2450 76680 2490
rect 76720 2450 76735 2490
rect 76665 2435 76735 2450
rect 77865 2490 77935 2520
rect 77865 2450 77880 2490
rect 77920 2450 77935 2490
rect 77865 2435 77935 2450
rect 8690 2250 8775 2265
rect 8690 2210 8705 2250
rect 8745 2210 8775 2250
rect 8690 2195 8775 2210
rect 10355 2250 10440 2265
rect 10355 2210 10385 2250
rect 10425 2210 10440 2250
rect 10355 2195 10440 2210
rect 13645 2250 13730 2265
rect 13645 2210 13660 2250
rect 13700 2210 13730 2250
rect 13645 2195 13730 2210
rect 15310 2250 15395 2265
rect 15310 2210 15340 2250
rect 15380 2210 15395 2250
rect 15310 2195 15395 2210
rect 18600 2250 18685 2265
rect 18600 2210 18615 2250
rect 18655 2210 18685 2250
rect 18600 2195 18685 2210
rect 20265 2250 20350 2265
rect 20265 2210 20295 2250
rect 20335 2210 20350 2250
rect 20265 2195 20350 2210
rect 23555 2250 23640 2265
rect 23555 2210 23570 2250
rect 23610 2210 23640 2250
rect 23555 2195 23640 2210
rect 25220 2250 25305 2265
rect 25220 2210 25250 2250
rect 25290 2210 25305 2250
rect 25220 2195 25305 2210
rect 28510 2250 28595 2265
rect 28510 2210 28525 2250
rect 28565 2210 28595 2250
rect 28510 2195 28595 2210
rect 30175 2250 30260 2265
rect 30175 2210 30205 2250
rect 30245 2210 30260 2250
rect 30175 2195 30260 2210
rect 33465 2250 33550 2265
rect 33465 2210 33480 2250
rect 33520 2210 33550 2250
rect 33465 2195 33550 2210
rect 35130 2250 35215 2265
rect 35130 2210 35160 2250
rect 35200 2210 35215 2250
rect 35130 2195 35215 2210
rect 38420 2250 38505 2265
rect 38420 2210 38435 2250
rect 38475 2210 38505 2250
rect 38420 2195 38505 2210
rect 40085 2250 40170 2265
rect 40085 2210 40115 2250
rect 40155 2210 40170 2250
rect 40085 2195 40170 2210
rect 43375 2250 43460 2265
rect 43375 2210 43390 2250
rect 43430 2210 43460 2250
rect 43375 2195 43460 2210
rect 45040 2250 45125 2265
rect 45040 2210 45070 2250
rect 45110 2210 45125 2250
rect 45040 2195 45125 2210
rect 48330 2250 48415 2265
rect 48330 2210 48345 2250
rect 48385 2210 48415 2250
rect 48330 2195 48415 2210
rect 49995 2250 50080 2265
rect 49995 2210 50025 2250
rect 50065 2210 50080 2250
rect 49995 2195 50080 2210
rect 53285 2250 53370 2265
rect 53285 2210 53300 2250
rect 53340 2210 53370 2250
rect 53285 2195 53370 2210
rect 54950 2250 55035 2265
rect 54950 2210 54980 2250
rect 55020 2210 55035 2250
rect 54950 2195 55035 2210
rect 58240 2250 58325 2265
rect 58240 2210 58255 2250
rect 58295 2210 58325 2250
rect 58240 2195 58325 2210
rect 59905 2250 59990 2265
rect 59905 2210 59935 2250
rect 59975 2210 59990 2250
rect 59905 2195 59990 2210
rect 63195 2250 63280 2265
rect 63195 2210 63210 2250
rect 63250 2210 63280 2250
rect 63195 2195 63280 2210
rect 64860 2250 64945 2265
rect 64860 2210 64890 2250
rect 64930 2210 64945 2250
rect 64860 2195 64945 2210
rect 68150 2250 68235 2265
rect 68150 2210 68165 2250
rect 68205 2210 68235 2250
rect 68150 2195 68235 2210
rect 69815 2250 69900 2265
rect 69815 2210 69845 2250
rect 69885 2210 69900 2250
rect 69815 2195 69900 2210
rect 73105 2250 73190 2265
rect 73105 2210 73120 2250
rect 73160 2210 73190 2250
rect 73105 2195 73190 2210
rect 74770 2250 74855 2265
rect 74770 2210 74800 2250
rect 74840 2210 74855 2250
rect 74770 2195 74855 2210
rect 8690 330 8775 345
rect 8690 290 8705 330
rect 8745 290 8775 330
rect 8690 275 8775 290
rect 10355 330 10440 345
rect 10355 290 10385 330
rect 10425 290 10440 330
rect 10355 275 10440 290
rect 13645 330 13730 345
rect 13645 290 13660 330
rect 13700 290 13730 330
rect 13645 275 13730 290
rect 15310 330 15395 345
rect 15310 290 15340 330
rect 15380 290 15395 330
rect 15310 275 15395 290
rect 18600 330 18685 345
rect 18600 290 18615 330
rect 18655 290 18685 330
rect 18600 275 18685 290
rect 20265 330 20350 345
rect 20265 290 20295 330
rect 20335 290 20350 330
rect 20265 275 20350 290
rect 23555 330 23640 345
rect 23555 290 23570 330
rect 23610 290 23640 330
rect 23555 275 23640 290
rect 25220 330 25305 345
rect 25220 290 25250 330
rect 25290 290 25305 330
rect 25220 275 25305 290
rect 28510 330 28595 345
rect 28510 290 28525 330
rect 28565 290 28595 330
rect 28510 275 28595 290
rect 30175 330 30260 345
rect 30175 290 30205 330
rect 30245 290 30260 330
rect 30175 275 30260 290
rect 33465 330 33550 345
rect 33465 290 33480 330
rect 33520 290 33550 330
rect 33465 275 33550 290
rect 35130 330 35215 345
rect 35130 290 35160 330
rect 35200 290 35215 330
rect 35130 275 35215 290
rect 38420 330 38505 345
rect 38420 290 38435 330
rect 38475 290 38505 330
rect 38420 275 38505 290
rect 40085 330 40170 345
rect 40085 290 40115 330
rect 40155 290 40170 330
rect 40085 275 40170 290
rect 43375 330 43460 345
rect 43375 290 43390 330
rect 43430 290 43460 330
rect 43375 275 43460 290
rect 45040 330 45125 345
rect 45040 290 45070 330
rect 45110 290 45125 330
rect 45040 275 45125 290
rect 48330 330 48415 345
rect 48330 290 48345 330
rect 48385 290 48415 330
rect 48330 275 48415 290
rect 49995 330 50080 345
rect 49995 290 50025 330
rect 50065 290 50080 330
rect 49995 275 50080 290
rect 53285 330 53370 345
rect 53285 290 53300 330
rect 53340 290 53370 330
rect 53285 275 53370 290
rect 54950 330 55035 345
rect 54950 290 54980 330
rect 55020 290 55035 330
rect 54950 275 55035 290
rect 58240 330 58325 345
rect 58240 290 58255 330
rect 58295 290 58325 330
rect 58240 275 58325 290
rect 59905 330 59990 345
rect 59905 290 59935 330
rect 59975 290 59990 330
rect 59905 275 59990 290
rect 63195 330 63280 345
rect 63195 290 63210 330
rect 63250 290 63280 330
rect 63195 275 63280 290
rect 64860 330 64945 345
rect 64860 290 64890 330
rect 64930 290 64945 330
rect 64860 275 64945 290
rect 68150 330 68235 345
rect 68150 290 68165 330
rect 68205 290 68235 330
rect 68150 275 68235 290
rect 69815 330 69900 345
rect 69815 290 69845 330
rect 69885 290 69900 330
rect 69815 275 69900 290
rect 73105 330 73190 345
rect 73105 290 73120 330
rect 73160 290 73190 330
rect 73105 275 73190 290
rect 74770 330 74855 345
rect 74770 290 74800 330
rect 74840 290 74855 330
rect 74770 275 74855 290
<< psubdiffcont >>
rect 8705 11435 8745 11475
rect 10385 11435 10425 11475
rect 13660 11435 13700 11475
rect 15340 11435 15380 11475
rect 18615 11435 18655 11475
rect 20295 11435 20335 11475
rect 23570 11435 23610 11475
rect 25250 11435 25290 11475
rect 28525 11435 28565 11475
rect 30205 11435 30245 11475
rect 33480 11435 33520 11475
rect 35160 11435 35200 11475
rect 38435 11435 38475 11475
rect 40115 11435 40155 11475
rect 43390 11435 43430 11475
rect 45070 11435 45110 11475
rect 48345 11435 48385 11475
rect 50025 11435 50065 11475
rect 53300 11435 53340 11475
rect 54980 11435 55020 11475
rect 58255 11435 58295 11475
rect 59935 11435 59975 11475
rect 63210 11435 63250 11475
rect 64890 11435 64930 11475
rect 68165 11435 68205 11475
rect 69845 11435 69885 11475
rect 73120 11435 73160 11475
rect 74800 11435 74840 11475
rect 8705 9515 8745 9555
rect 10385 9515 10425 9555
rect 13660 9515 13700 9555
rect 15340 9515 15380 9555
rect 18615 9515 18655 9555
rect 20295 9515 20335 9555
rect 23570 9515 23610 9555
rect 25250 9515 25290 9555
rect 28525 9515 28565 9555
rect 30205 9515 30245 9555
rect 33480 9515 33520 9555
rect 35160 9515 35200 9555
rect 38435 9515 38475 9555
rect 40115 9515 40155 9555
rect 43390 9515 43430 9555
rect 45070 9515 45110 9555
rect 48345 9515 48385 9555
rect 50025 9515 50065 9555
rect 53300 9515 53340 9555
rect 54980 9515 55020 9555
rect 58255 9515 58295 9555
rect 59935 9515 59975 9555
rect 63210 9515 63250 9555
rect 64890 9515 64930 9555
rect 68165 9515 68205 9555
rect 69845 9515 69885 9555
rect 73120 9515 73160 9555
rect 74800 9515 74840 9555
rect 5630 9230 5670 9270
rect 6830 9230 6870 9270
rect 7310 9230 7350 9270
rect 8510 9230 8550 9270
rect 10585 9230 10625 9270
rect 11785 9230 11825 9270
rect 12265 9230 12305 9270
rect 13465 9230 13505 9270
rect 15540 9230 15580 9270
rect 16740 9230 16780 9270
rect 17220 9230 17260 9270
rect 18420 9230 18460 9270
rect 20495 9230 20535 9270
rect 21695 9230 21735 9270
rect 22175 9230 22215 9270
rect 23375 9230 23415 9270
rect 25450 9230 25490 9270
rect 26650 9230 26690 9270
rect 27130 9230 27170 9270
rect 28330 9230 28370 9270
rect 30405 9230 30445 9270
rect 31605 9230 31645 9270
rect 32085 9230 32125 9270
rect 33285 9230 33325 9270
rect 35360 9230 35400 9270
rect 36560 9230 36600 9270
rect 37040 9230 37080 9270
rect 38240 9230 38280 9270
rect 40315 9230 40355 9270
rect 41515 9230 41555 9270
rect 41995 9230 42035 9270
rect 43195 9230 43235 9270
rect 45270 9230 45310 9270
rect 46470 9230 46510 9270
rect 46950 9230 46990 9270
rect 48150 9230 48190 9270
rect 50225 9230 50265 9270
rect 51425 9230 51465 9270
rect 51905 9230 51945 9270
rect 53105 9230 53145 9270
rect 55180 9230 55220 9270
rect 56380 9230 56420 9270
rect 56860 9230 56900 9270
rect 58060 9230 58100 9270
rect 60135 9230 60175 9270
rect 61335 9230 61375 9270
rect 61815 9230 61855 9270
rect 63015 9230 63055 9270
rect 65090 9230 65130 9270
rect 66290 9230 66330 9270
rect 66770 9230 66810 9270
rect 67970 9230 68010 9270
rect 70045 9230 70085 9270
rect 71245 9230 71285 9270
rect 71725 9230 71765 9270
rect 72925 9230 72965 9270
rect 75000 9230 75040 9270
rect 76200 9230 76240 9270
rect 76680 9230 76720 9270
rect 77880 9230 77920 9270
rect 5630 8600 5670 8640
rect 6830 8600 6870 8640
rect 7310 8600 7350 8640
rect 8510 8600 8550 8640
rect 10585 8600 10625 8640
rect 11785 8600 11825 8640
rect 12265 8600 12305 8640
rect 13465 8600 13505 8640
rect 15540 8600 15580 8640
rect 16740 8600 16780 8640
rect 17220 8600 17260 8640
rect 18420 8600 18460 8640
rect 20495 8600 20535 8640
rect 21695 8600 21735 8640
rect 22175 8600 22215 8640
rect 23375 8600 23415 8640
rect 25450 8600 25490 8640
rect 26650 8600 26690 8640
rect 27130 8600 27170 8640
rect 28330 8600 28370 8640
rect 30405 8600 30445 8640
rect 31605 8600 31645 8640
rect 32085 8600 32125 8640
rect 33285 8600 33325 8640
rect 35360 8600 35400 8640
rect 36560 8600 36600 8640
rect 37040 8600 37080 8640
rect 38240 8600 38280 8640
rect 40315 8600 40355 8640
rect 41515 8600 41555 8640
rect 41995 8600 42035 8640
rect 43195 8600 43235 8640
rect 45270 8600 45310 8640
rect 46470 8600 46510 8640
rect 46950 8600 46990 8640
rect 48150 8600 48190 8640
rect 50225 8600 50265 8640
rect 51425 8600 51465 8640
rect 51905 8600 51945 8640
rect 53105 8600 53145 8640
rect 55180 8600 55220 8640
rect 56380 8600 56420 8640
rect 56860 8600 56900 8640
rect 58060 8600 58100 8640
rect 60135 8600 60175 8640
rect 61335 8600 61375 8640
rect 61815 8600 61855 8640
rect 63015 8600 63055 8640
rect 65090 8600 65130 8640
rect 66290 8600 66330 8640
rect 66770 8600 66810 8640
rect 67970 8600 68010 8640
rect 70045 8600 70085 8640
rect 71245 8600 71285 8640
rect 71725 8600 71765 8640
rect 72925 8600 72965 8640
rect 75000 8600 75040 8640
rect 76200 8600 76240 8640
rect 76680 8600 76720 8640
rect 77880 8600 77920 8640
rect 8705 8360 8745 8400
rect 10385 8360 10425 8400
rect 13660 8360 13700 8400
rect 15340 8360 15380 8400
rect 18615 8360 18655 8400
rect 20295 8360 20335 8400
rect 23570 8360 23610 8400
rect 25250 8360 25290 8400
rect 28525 8360 28565 8400
rect 30205 8360 30245 8400
rect 33480 8360 33520 8400
rect 35160 8360 35200 8400
rect 38435 8360 38475 8400
rect 40115 8360 40155 8400
rect 43390 8360 43430 8400
rect 45070 8360 45110 8400
rect 48345 8360 48385 8400
rect 50025 8360 50065 8400
rect 53300 8360 53340 8400
rect 54980 8360 55020 8400
rect 58255 8360 58295 8400
rect 59935 8360 59975 8400
rect 63210 8360 63250 8400
rect 64890 8360 64930 8400
rect 68165 8360 68205 8400
rect 69845 8360 69885 8400
rect 73120 8360 73160 8400
rect 74800 8360 74840 8400
rect 8705 6440 8745 6480
rect 10385 6440 10425 6480
rect 13660 6440 13700 6480
rect 15340 6440 15380 6480
rect 18615 6440 18655 6480
rect 20295 6440 20335 6480
rect 23570 6440 23610 6480
rect 25250 6440 25290 6480
rect 28525 6440 28565 6480
rect 30205 6440 30245 6480
rect 33480 6440 33520 6480
rect 35160 6440 35200 6480
rect 38435 6440 38475 6480
rect 40115 6440 40155 6480
rect 43390 6440 43430 6480
rect 45070 6440 45110 6480
rect 48345 6440 48385 6480
rect 50025 6440 50065 6480
rect 53300 6440 53340 6480
rect 54980 6440 55020 6480
rect 58255 6440 58295 6480
rect 59935 6440 59975 6480
rect 63210 6440 63250 6480
rect 64890 6440 64930 6480
rect 68165 6440 68205 6480
rect 69845 6440 69885 6480
rect 73120 6440 73160 6480
rect 74800 6440 74840 6480
rect 5630 6155 5670 6195
rect 6830 6155 6870 6195
rect 7310 6155 7350 6195
rect 8510 6155 8550 6195
rect 10585 6155 10625 6195
rect 11785 6155 11825 6195
rect 12265 6155 12305 6195
rect 13465 6155 13505 6195
rect 15540 6155 15580 6195
rect 16740 6155 16780 6195
rect 17220 6155 17260 6195
rect 18420 6155 18460 6195
rect 20495 6155 20535 6195
rect 21695 6155 21735 6195
rect 22175 6155 22215 6195
rect 23375 6155 23415 6195
rect 25450 6155 25490 6195
rect 26650 6155 26690 6195
rect 27130 6155 27170 6195
rect 28330 6155 28370 6195
rect 30405 6155 30445 6195
rect 31605 6155 31645 6195
rect 32085 6155 32125 6195
rect 33285 6155 33325 6195
rect 35360 6155 35400 6195
rect 36560 6155 36600 6195
rect 37040 6155 37080 6195
rect 38240 6155 38280 6195
rect 40315 6155 40355 6195
rect 41515 6155 41555 6195
rect 41995 6155 42035 6195
rect 43195 6155 43235 6195
rect 45270 6155 45310 6195
rect 46470 6155 46510 6195
rect 46950 6155 46990 6195
rect 48150 6155 48190 6195
rect 50225 6155 50265 6195
rect 51425 6155 51465 6195
rect 51905 6155 51945 6195
rect 53105 6155 53145 6195
rect 55180 6155 55220 6195
rect 56380 6155 56420 6195
rect 56860 6155 56900 6195
rect 58060 6155 58100 6195
rect 60135 6155 60175 6195
rect 61335 6155 61375 6195
rect 61815 6155 61855 6195
rect 63015 6155 63055 6195
rect 65090 6155 65130 6195
rect 66290 6155 66330 6195
rect 66770 6155 66810 6195
rect 67970 6155 68010 6195
rect 70045 6155 70085 6195
rect 71245 6155 71285 6195
rect 71725 6155 71765 6195
rect 72925 6155 72965 6195
rect 75000 6155 75040 6195
rect 76200 6155 76240 6195
rect 76680 6155 76720 6195
rect 77880 6155 77920 6195
rect 5630 5525 5670 5565
rect 6830 5525 6870 5565
rect 7310 5525 7350 5565
rect 8510 5525 8550 5565
rect 10585 5525 10625 5565
rect 11785 5525 11825 5565
rect 12265 5525 12305 5565
rect 13465 5525 13505 5565
rect 15540 5525 15580 5565
rect 16740 5525 16780 5565
rect 17220 5525 17260 5565
rect 18420 5525 18460 5565
rect 20495 5525 20535 5565
rect 21695 5525 21735 5565
rect 22175 5525 22215 5565
rect 23375 5525 23415 5565
rect 25450 5525 25490 5565
rect 26650 5525 26690 5565
rect 27130 5525 27170 5565
rect 28330 5525 28370 5565
rect 30405 5525 30445 5565
rect 31605 5525 31645 5565
rect 32085 5525 32125 5565
rect 33285 5525 33325 5565
rect 35360 5525 35400 5565
rect 36560 5525 36600 5565
rect 37040 5525 37080 5565
rect 38240 5525 38280 5565
rect 40315 5525 40355 5565
rect 41515 5525 41555 5565
rect 41995 5525 42035 5565
rect 43195 5525 43235 5565
rect 45270 5525 45310 5565
rect 46470 5525 46510 5565
rect 46950 5525 46990 5565
rect 48150 5525 48190 5565
rect 50225 5525 50265 5565
rect 51425 5525 51465 5565
rect 51905 5525 51945 5565
rect 53105 5525 53145 5565
rect 55180 5525 55220 5565
rect 56380 5525 56420 5565
rect 56860 5525 56900 5565
rect 58060 5525 58100 5565
rect 60135 5525 60175 5565
rect 61335 5525 61375 5565
rect 61815 5525 61855 5565
rect 63015 5525 63055 5565
rect 65090 5525 65130 5565
rect 66290 5525 66330 5565
rect 66770 5525 66810 5565
rect 67970 5525 68010 5565
rect 70045 5525 70085 5565
rect 71245 5525 71285 5565
rect 71725 5525 71765 5565
rect 72925 5525 72965 5565
rect 75000 5525 75040 5565
rect 76200 5525 76240 5565
rect 76680 5525 76720 5565
rect 77880 5525 77920 5565
rect 8705 5285 8745 5325
rect 10385 5285 10425 5325
rect 13660 5285 13700 5325
rect 15340 5285 15380 5325
rect 18615 5285 18655 5325
rect 20295 5285 20335 5325
rect 23570 5285 23610 5325
rect 25250 5285 25290 5325
rect 28525 5285 28565 5325
rect 30205 5285 30245 5325
rect 33480 5285 33520 5325
rect 35160 5285 35200 5325
rect 38435 5285 38475 5325
rect 40115 5285 40155 5325
rect 43390 5285 43430 5325
rect 45070 5285 45110 5325
rect 48345 5285 48385 5325
rect 50025 5285 50065 5325
rect 53300 5285 53340 5325
rect 54980 5285 55020 5325
rect 58255 5285 58295 5325
rect 59935 5285 59975 5325
rect 63210 5285 63250 5325
rect 64890 5285 64930 5325
rect 68165 5285 68205 5325
rect 69845 5285 69885 5325
rect 73120 5285 73160 5325
rect 74800 5285 74840 5325
rect 8705 3365 8745 3405
rect 10385 3365 10425 3405
rect 13660 3365 13700 3405
rect 15340 3365 15380 3405
rect 18615 3365 18655 3405
rect 20295 3365 20335 3405
rect 23570 3365 23610 3405
rect 25250 3365 25290 3405
rect 28525 3365 28565 3405
rect 30205 3365 30245 3405
rect 33480 3365 33520 3405
rect 35160 3365 35200 3405
rect 38435 3365 38475 3405
rect 40115 3365 40155 3405
rect 43390 3365 43430 3405
rect 45070 3365 45110 3405
rect 48345 3365 48385 3405
rect 50025 3365 50065 3405
rect 53300 3365 53340 3405
rect 54980 3365 55020 3405
rect 58255 3365 58295 3405
rect 59935 3365 59975 3405
rect 63210 3365 63250 3405
rect 64890 3365 64930 3405
rect 68165 3365 68205 3405
rect 69845 3365 69885 3405
rect 73120 3365 73160 3405
rect 74800 3365 74840 3405
rect 675 3080 715 3120
rect 5630 3080 5670 3120
rect 6830 3080 6870 3120
rect 7310 3080 7350 3120
rect 8510 3080 8550 3120
rect 10585 3080 10625 3120
rect 11785 3080 11825 3120
rect 12265 3080 12305 3120
rect 13465 3080 13505 3120
rect 15540 3080 15580 3120
rect 16740 3080 16780 3120
rect 17220 3080 17260 3120
rect 18420 3080 18460 3120
rect 20495 3080 20535 3120
rect 21695 3080 21735 3120
rect 22175 3080 22215 3120
rect 23375 3080 23415 3120
rect 25450 3080 25490 3120
rect 26650 3080 26690 3120
rect 27130 3080 27170 3120
rect 28330 3080 28370 3120
rect 30405 3080 30445 3120
rect 31605 3080 31645 3120
rect 32085 3080 32125 3120
rect 33285 3080 33325 3120
rect 35360 3080 35400 3120
rect 36560 3080 36600 3120
rect 37040 3080 37080 3120
rect 38240 3080 38280 3120
rect 40315 3080 40355 3120
rect 41515 3080 41555 3120
rect 41995 3080 42035 3120
rect 43195 3080 43235 3120
rect 45270 3080 45310 3120
rect 46470 3080 46510 3120
rect 46950 3080 46990 3120
rect 48150 3080 48190 3120
rect 50225 3080 50265 3120
rect 51425 3080 51465 3120
rect 51905 3080 51945 3120
rect 53105 3080 53145 3120
rect 55180 3080 55220 3120
rect 56380 3080 56420 3120
rect 56860 3080 56900 3120
rect 58060 3080 58100 3120
rect 60135 3080 60175 3120
rect 61335 3080 61375 3120
rect 61815 3080 61855 3120
rect 63015 3080 63055 3120
rect 65090 3080 65130 3120
rect 66290 3080 66330 3120
rect 66770 3080 66810 3120
rect 67970 3080 68010 3120
rect 70045 3080 70085 3120
rect 71245 3080 71285 3120
rect 71725 3080 71765 3120
rect 72925 3080 72965 3120
rect 75000 3080 75040 3120
rect 76200 3080 76240 3120
rect 76680 3080 76720 3120
rect 77880 3080 77920 3120
rect 675 2450 715 2490
rect 5630 2450 5670 2490
rect 6830 2450 6870 2490
rect 7310 2450 7350 2490
rect 8510 2450 8550 2490
rect 10585 2450 10625 2490
rect 11785 2450 11825 2490
rect 12265 2450 12305 2490
rect 13465 2450 13505 2490
rect 15540 2450 15580 2490
rect 16740 2450 16780 2490
rect 17220 2450 17260 2490
rect 18420 2450 18460 2490
rect 20495 2450 20535 2490
rect 21695 2450 21735 2490
rect 22175 2450 22215 2490
rect 23375 2450 23415 2490
rect 25450 2450 25490 2490
rect 26650 2450 26690 2490
rect 27130 2450 27170 2490
rect 28330 2450 28370 2490
rect 30405 2450 30445 2490
rect 31605 2450 31645 2490
rect 32085 2450 32125 2490
rect 33285 2450 33325 2490
rect 35360 2450 35400 2490
rect 36560 2450 36600 2490
rect 37040 2450 37080 2490
rect 38240 2450 38280 2490
rect 40315 2450 40355 2490
rect 41515 2450 41555 2490
rect 41995 2450 42035 2490
rect 43195 2450 43235 2490
rect 45270 2450 45310 2490
rect 46470 2450 46510 2490
rect 46950 2450 46990 2490
rect 48150 2450 48190 2490
rect 50225 2450 50265 2490
rect 51425 2450 51465 2490
rect 51905 2450 51945 2490
rect 53105 2450 53145 2490
rect 55180 2450 55220 2490
rect 56380 2450 56420 2490
rect 56860 2450 56900 2490
rect 58060 2450 58100 2490
rect 60135 2450 60175 2490
rect 61335 2450 61375 2490
rect 61815 2450 61855 2490
rect 63015 2450 63055 2490
rect 65090 2450 65130 2490
rect 66290 2450 66330 2490
rect 66770 2450 66810 2490
rect 67970 2450 68010 2490
rect 70045 2450 70085 2490
rect 71245 2450 71285 2490
rect 71725 2450 71765 2490
rect 72925 2450 72965 2490
rect 75000 2450 75040 2490
rect 76200 2450 76240 2490
rect 76680 2450 76720 2490
rect 77880 2450 77920 2490
rect 8705 2210 8745 2250
rect 10385 2210 10425 2250
rect 13660 2210 13700 2250
rect 15340 2210 15380 2250
rect 18615 2210 18655 2250
rect 20295 2210 20335 2250
rect 23570 2210 23610 2250
rect 25250 2210 25290 2250
rect 28525 2210 28565 2250
rect 30205 2210 30245 2250
rect 33480 2210 33520 2250
rect 35160 2210 35200 2250
rect 38435 2210 38475 2250
rect 40115 2210 40155 2250
rect 43390 2210 43430 2250
rect 45070 2210 45110 2250
rect 48345 2210 48385 2250
rect 50025 2210 50065 2250
rect 53300 2210 53340 2250
rect 54980 2210 55020 2250
rect 58255 2210 58295 2250
rect 59935 2210 59975 2250
rect 63210 2210 63250 2250
rect 64890 2210 64930 2250
rect 68165 2210 68205 2250
rect 69845 2210 69885 2250
rect 73120 2210 73160 2250
rect 74800 2210 74840 2250
rect 8705 290 8745 330
rect 10385 290 10425 330
rect 13660 290 13700 330
rect 15340 290 15380 330
rect 18615 290 18655 330
rect 20295 290 20335 330
rect 23570 290 23610 330
rect 25250 290 25290 330
rect 28525 290 28565 330
rect 30205 290 30245 330
rect 33480 290 33520 330
rect 35160 290 35200 330
rect 38435 290 38475 330
rect 40115 290 40155 330
rect 43390 290 43430 330
rect 45070 290 45110 330
rect 48345 290 48385 330
rect 50025 290 50065 330
rect 53300 290 53340 330
rect 54980 290 55020 330
rect 58255 290 58295 330
rect 59935 290 59975 330
rect 63210 290 63250 330
rect 64890 290 64930 330
rect 68165 290 68205 330
rect 69845 290 69885 330
rect 73120 290 73160 330
rect 74800 290 74840 330
<< poly >>
rect 7045 40 7130 55
rect 7045 -10 7060 40
rect 7115 -10 7130 40
rect 7045 -25 7130 -10
rect 12000 40 12085 55
rect 12000 -10 12015 40
rect 12070 -10 12085 40
rect 12000 -25 12085 -10
rect 16955 40 17040 55
rect 16955 -10 16970 40
rect 17025 -10 17040 40
rect 16955 -25 17040 -10
rect 21910 40 21995 55
rect 21910 -10 21925 40
rect 21980 -10 21995 40
rect 21910 -25 21995 -10
rect 26865 40 26950 55
rect 26865 -10 26880 40
rect 26935 -10 26950 40
rect 26865 -25 26950 -10
rect 31820 40 31905 55
rect 31820 -10 31835 40
rect 31890 -10 31905 40
rect 31820 -25 31905 -10
rect 36775 40 36860 55
rect 36775 -10 36790 40
rect 36845 -10 36860 40
rect 36775 -25 36860 -10
rect 41730 40 41815 55
rect 41730 -10 41745 40
rect 41800 -10 41815 40
rect 41730 -25 41815 -10
rect 46685 40 46770 55
rect 46685 -10 46700 40
rect 46755 -10 46770 40
rect 46685 -25 46770 -10
rect 51640 40 51725 55
rect 51640 -10 51655 40
rect 51710 -10 51725 40
rect 51640 -25 51725 -10
rect 56595 40 56680 55
rect 56595 -10 56610 40
rect 56665 -10 56680 40
rect 56595 -25 56680 -10
rect 61550 40 61635 55
rect 61550 -10 61565 40
rect 61620 -10 61635 40
rect 61550 -25 61635 -10
rect 66505 40 66590 55
rect 66505 -10 66520 40
rect 66575 -10 66590 40
rect 66505 -25 66590 -10
rect 71460 40 71545 55
rect 71460 -10 71475 40
rect 71530 -10 71545 40
rect 71460 -25 71545 -10
rect 76415 40 76500 55
rect 76415 -10 76430 40
rect 76485 -10 76500 40
rect 76415 -25 76500 -10
<< polycont >>
rect 7060 -10 7115 40
rect 12015 -10 12070 40
rect 16970 -10 17025 40
rect 21925 -10 21980 40
rect 26880 -10 26935 40
rect 31835 -10 31890 40
rect 36790 -10 36845 40
rect 41745 -10 41800 40
rect 46700 -10 46755 40
rect 51655 -10 51710 40
rect 56610 -10 56665 40
rect 61565 -10 61620 40
rect 66520 -10 66575 40
rect 71475 -10 71530 40
rect 76430 -10 76485 40
<< locali >>
rect -345 12050 78830 12065
rect -345 11920 -330 12050
rect -200 11985 78830 12050
rect -200 11920 -185 11985
rect -345 11905 -185 11920
rect 2090 11745 2175 11985
rect 7045 11745 7130 11985
rect 12000 11745 12085 11985
rect 16955 11745 17040 11985
rect 21910 11745 21995 11985
rect 26865 11745 26950 11985
rect 31820 11745 31905 11985
rect 36775 11745 36860 11985
rect 41730 11745 41815 11985
rect 46685 11745 46770 11985
rect 51640 11745 51725 11985
rect 56595 11745 56680 11985
rect 61550 11745 61635 11985
rect 66505 11745 66590 11985
rect 71460 11745 71545 11985
rect 76415 11745 76500 11985
rect 3735 11420 5485 11490
rect 8690 11475 10440 11490
rect 8690 11435 8705 11475
rect 8745 11435 10385 11475
rect 10425 11435 10440 11475
rect 8690 11420 10440 11435
rect 13645 11475 15395 11490
rect 13645 11435 13660 11475
rect 13700 11435 15340 11475
rect 15380 11435 15395 11475
rect 13645 11420 15395 11435
rect 18600 11475 20350 11490
rect 18600 11435 18615 11475
rect 18655 11435 20295 11475
rect 20335 11435 20350 11475
rect 18600 11420 20350 11435
rect 23555 11475 25305 11490
rect 23555 11435 23570 11475
rect 23610 11435 25250 11475
rect 25290 11435 25305 11475
rect 23555 11420 25305 11435
rect 28510 11475 30260 11490
rect 28510 11435 28525 11475
rect 28565 11435 30205 11475
rect 30245 11435 30260 11475
rect 28510 11420 30260 11435
rect 33465 11475 35215 11490
rect 33465 11435 33480 11475
rect 33520 11435 35160 11475
rect 35200 11435 35215 11475
rect 33465 11420 35215 11435
rect 38420 11475 40170 11490
rect 38420 11435 38435 11475
rect 38475 11435 40115 11475
rect 40155 11435 40170 11475
rect 38420 11420 40170 11435
rect 43375 11475 45125 11490
rect 43375 11435 43390 11475
rect 43430 11435 45070 11475
rect 45110 11435 45125 11475
rect 43375 11420 45125 11435
rect 48330 11475 50080 11490
rect 48330 11435 48345 11475
rect 48385 11435 50025 11475
rect 50065 11435 50080 11475
rect 48330 11420 50080 11435
rect 53285 11475 55035 11490
rect 53285 11435 53300 11475
rect 53340 11435 54980 11475
rect 55020 11435 55035 11475
rect 53285 11420 55035 11435
rect 58240 11475 59990 11490
rect 58240 11435 58255 11475
rect 58295 11435 59935 11475
rect 59975 11435 59990 11475
rect 58240 11420 59990 11435
rect 63195 11475 64945 11490
rect 63195 11435 63210 11475
rect 63250 11435 64890 11475
rect 64930 11435 64945 11475
rect 63195 11420 64945 11435
rect 68150 11475 69900 11490
rect 68150 11435 68165 11475
rect 68205 11435 69845 11475
rect 69885 11435 69900 11475
rect 68150 11420 69900 11435
rect 73105 11475 74855 11490
rect 73105 11435 73120 11475
rect 73160 11435 74800 11475
rect 74840 11435 74855 11475
rect 73105 11420 74855 11435
rect 4595 9570 4670 11420
rect 9550 9570 9625 11420
rect 14505 9570 14580 11420
rect 19460 9570 19535 11420
rect 24415 9570 24490 11420
rect 29370 9570 29445 11420
rect 34325 9570 34400 11420
rect 39280 9570 39355 11420
rect 44235 9570 44310 11420
rect 49190 9570 49265 11420
rect 54145 9570 54220 11420
rect 59100 9570 59175 11420
rect 64055 9570 64130 11420
rect 69010 9570 69085 11420
rect 73965 9570 74040 11420
rect 3735 9500 5485 9570
rect 8690 9555 10440 9570
rect 8690 9515 8705 9555
rect 8745 9515 10385 9555
rect 10425 9515 10440 9555
rect 8690 9500 10440 9515
rect 13645 9555 15395 9570
rect 13645 9515 13660 9555
rect 13700 9515 15340 9555
rect 15380 9515 15395 9555
rect 13645 9500 15395 9515
rect 18600 9555 20350 9570
rect 18600 9515 18615 9555
rect 18655 9515 20295 9555
rect 20335 9515 20350 9555
rect 18600 9500 20350 9515
rect 23555 9555 25305 9570
rect 23555 9515 23570 9555
rect 23610 9515 25250 9555
rect 25290 9515 25305 9555
rect 23555 9500 25305 9515
rect 28510 9555 30260 9570
rect 28510 9515 28525 9555
rect 28565 9515 30205 9555
rect 30245 9515 30260 9555
rect 28510 9500 30260 9515
rect 33465 9555 35215 9570
rect 33465 9515 33480 9555
rect 33520 9515 35160 9555
rect 35200 9515 35215 9555
rect 33465 9500 35215 9515
rect 38420 9555 40170 9570
rect 38420 9515 38435 9555
rect 38475 9515 40115 9555
rect 40155 9515 40170 9555
rect 38420 9500 40170 9515
rect 43375 9555 45125 9570
rect 43375 9515 43390 9555
rect 43430 9515 45070 9555
rect 45110 9515 45125 9555
rect 43375 9500 45125 9515
rect 48330 9555 50080 9570
rect 48330 9515 48345 9555
rect 48385 9515 50025 9555
rect 50065 9515 50080 9555
rect 48330 9500 50080 9515
rect 53285 9555 55035 9570
rect 53285 9515 53300 9555
rect 53340 9515 54980 9555
rect 55020 9515 55035 9555
rect 53285 9500 55035 9515
rect 58240 9555 59990 9570
rect 58240 9515 58255 9555
rect 58295 9515 59935 9555
rect 59975 9515 59990 9555
rect 58240 9500 59990 9515
rect 63195 9555 64945 9570
rect 63195 9515 63210 9555
rect 63250 9515 64890 9555
rect 64930 9515 64945 9555
rect 63195 9500 64945 9515
rect 68150 9555 69900 9570
rect 68150 9515 68165 9555
rect 68205 9515 69845 9555
rect 69885 9515 69900 9555
rect 68150 9500 69900 9515
rect 73105 9555 74855 9570
rect 73105 9515 73120 9555
rect 73160 9515 74800 9555
rect 74840 9515 74855 9555
rect 73105 9500 74855 9515
rect 660 8935 730 9285
rect 660 8900 675 8935
rect 715 8900 730 8935
rect 660 8585 730 8900
rect 1860 8935 1930 9285
rect 1860 8900 1875 8935
rect 1915 8900 1930 8935
rect 1860 8585 1930 8900
rect 2090 8670 2175 9200
rect 2340 8935 2410 9285
rect 2340 8900 2355 8935
rect 2395 8900 2410 8935
rect 2340 8585 2410 8900
rect 3540 8935 3610 9285
rect 3540 8900 3555 8935
rect 3595 8900 3610 8935
rect 3540 8585 3610 8900
rect 4595 8415 4670 9500
rect 5615 9270 5685 9285
rect 5615 9230 5630 9270
rect 5670 9230 5685 9270
rect 5615 8935 5685 9230
rect 5615 8900 5630 8935
rect 5670 8900 5685 8935
rect 5615 8640 5685 8900
rect 5615 8600 5630 8640
rect 5670 8600 5685 8640
rect 5615 8585 5685 8600
rect 6815 9270 6885 9285
rect 6815 9230 6830 9270
rect 6870 9230 6885 9270
rect 6815 8935 6885 9230
rect 7295 9270 7365 9285
rect 7295 9230 7310 9270
rect 7350 9230 7365 9270
rect 6815 8900 6830 8935
rect 6870 8900 6885 8935
rect 6815 8640 6885 8900
rect 7045 8670 7130 9200
rect 7295 8935 7365 9230
rect 7295 8900 7310 8935
rect 7350 8900 7365 8935
rect 6815 8600 6830 8640
rect 6870 8600 6885 8640
rect 6815 8585 6885 8600
rect 7295 8640 7365 8900
rect 7295 8600 7310 8640
rect 7350 8600 7365 8640
rect 7295 8585 7365 8600
rect 8495 9270 8565 9285
rect 8495 9230 8510 9270
rect 8550 9230 8565 9270
rect 8495 8935 8565 9230
rect 8495 8900 8510 8935
rect 8550 8900 8565 8935
rect 8495 8640 8565 8900
rect 8495 8600 8510 8640
rect 8550 8600 8565 8640
rect 8495 8585 8565 8600
rect 9550 8415 9625 9500
rect 10570 9270 10640 9285
rect 10570 9230 10585 9270
rect 10625 9230 10640 9270
rect 10570 8935 10640 9230
rect 10570 8900 10585 8935
rect 10625 8900 10640 8935
rect 10570 8640 10640 8900
rect 10570 8600 10585 8640
rect 10625 8600 10640 8640
rect 10570 8585 10640 8600
rect 11770 9270 11840 9285
rect 11770 9230 11785 9270
rect 11825 9230 11840 9270
rect 11770 8935 11840 9230
rect 12250 9270 12320 9285
rect 12250 9230 12265 9270
rect 12305 9230 12320 9270
rect 11770 8900 11785 8935
rect 11825 8900 11840 8935
rect 11770 8640 11840 8900
rect 12000 8670 12085 9200
rect 12250 8935 12320 9230
rect 12250 8900 12265 8935
rect 12305 8900 12320 8935
rect 11770 8600 11785 8640
rect 11825 8600 11840 8640
rect 11770 8585 11840 8600
rect 12250 8640 12320 8900
rect 12250 8600 12265 8640
rect 12305 8600 12320 8640
rect 12250 8585 12320 8600
rect 13450 9270 13520 9285
rect 13450 9230 13465 9270
rect 13505 9230 13520 9270
rect 13450 8935 13520 9230
rect 13450 8900 13465 8935
rect 13505 8900 13520 8935
rect 13450 8640 13520 8900
rect 13450 8600 13465 8640
rect 13505 8600 13520 8640
rect 13450 8585 13520 8600
rect 14505 8415 14580 9500
rect 15525 9270 15595 9285
rect 15525 9230 15540 9270
rect 15580 9230 15595 9270
rect 15525 8935 15595 9230
rect 15525 8900 15540 8935
rect 15580 8900 15595 8935
rect 15525 8640 15595 8900
rect 15525 8600 15540 8640
rect 15580 8600 15595 8640
rect 15525 8585 15595 8600
rect 16725 9270 16795 9285
rect 16725 9230 16740 9270
rect 16780 9230 16795 9270
rect 16725 8935 16795 9230
rect 17205 9270 17275 9285
rect 17205 9230 17220 9270
rect 17260 9230 17275 9270
rect 16725 8900 16740 8935
rect 16780 8900 16795 8935
rect 16725 8640 16795 8900
rect 16955 8670 17040 9200
rect 17205 8935 17275 9230
rect 17205 8900 17220 8935
rect 17260 8900 17275 8935
rect 16725 8600 16740 8640
rect 16780 8600 16795 8640
rect 16725 8585 16795 8600
rect 17205 8640 17275 8900
rect 17205 8600 17220 8640
rect 17260 8600 17275 8640
rect 17205 8585 17275 8600
rect 18405 9270 18475 9285
rect 18405 9230 18420 9270
rect 18460 9230 18475 9270
rect 18405 8935 18475 9230
rect 18405 8900 18420 8935
rect 18460 8900 18475 8935
rect 18405 8640 18475 8900
rect 18405 8600 18420 8640
rect 18460 8600 18475 8640
rect 18405 8585 18475 8600
rect 19460 8415 19535 9500
rect 20480 9270 20550 9285
rect 20480 9230 20495 9270
rect 20535 9230 20550 9270
rect 20480 8935 20550 9230
rect 20480 8900 20495 8935
rect 20535 8900 20550 8935
rect 20480 8640 20550 8900
rect 20480 8600 20495 8640
rect 20535 8600 20550 8640
rect 20480 8585 20550 8600
rect 21680 9270 21750 9285
rect 21680 9230 21695 9270
rect 21735 9230 21750 9270
rect 21680 8935 21750 9230
rect 22160 9270 22230 9285
rect 22160 9230 22175 9270
rect 22215 9230 22230 9270
rect 21680 8900 21695 8935
rect 21735 8900 21750 8935
rect 21680 8640 21750 8900
rect 21910 8670 21995 9200
rect 22160 8935 22230 9230
rect 22160 8900 22175 8935
rect 22215 8900 22230 8935
rect 21680 8600 21695 8640
rect 21735 8600 21750 8640
rect 21680 8585 21750 8600
rect 22160 8640 22230 8900
rect 22160 8600 22175 8640
rect 22215 8600 22230 8640
rect 22160 8585 22230 8600
rect 23360 9270 23430 9285
rect 23360 9230 23375 9270
rect 23415 9230 23430 9270
rect 23360 8935 23430 9230
rect 23360 8900 23375 8935
rect 23415 8900 23430 8935
rect 23360 8640 23430 8900
rect 23360 8600 23375 8640
rect 23415 8600 23430 8640
rect 23360 8585 23430 8600
rect 24415 8415 24490 9500
rect 25435 9270 25505 9285
rect 25435 9230 25450 9270
rect 25490 9230 25505 9270
rect 25435 8935 25505 9230
rect 25435 8900 25450 8935
rect 25490 8900 25505 8935
rect 25435 8640 25505 8900
rect 25435 8600 25450 8640
rect 25490 8600 25505 8640
rect 25435 8585 25505 8600
rect 26635 9270 26705 9285
rect 26635 9230 26650 9270
rect 26690 9230 26705 9270
rect 26635 8935 26705 9230
rect 27115 9270 27185 9285
rect 27115 9230 27130 9270
rect 27170 9230 27185 9270
rect 26635 8900 26650 8935
rect 26690 8900 26705 8935
rect 26635 8640 26705 8900
rect 26865 8670 26950 9200
rect 27115 8935 27185 9230
rect 27115 8900 27130 8935
rect 27170 8900 27185 8935
rect 26635 8600 26650 8640
rect 26690 8600 26705 8640
rect 26635 8585 26705 8600
rect 27115 8640 27185 8900
rect 27115 8600 27130 8640
rect 27170 8600 27185 8640
rect 27115 8585 27185 8600
rect 28315 9270 28385 9285
rect 28315 9230 28330 9270
rect 28370 9230 28385 9270
rect 28315 8935 28385 9230
rect 28315 8900 28330 8935
rect 28370 8900 28385 8935
rect 28315 8640 28385 8900
rect 28315 8600 28330 8640
rect 28370 8600 28385 8640
rect 28315 8585 28385 8600
rect 29370 8415 29445 9500
rect 30390 9270 30460 9285
rect 30390 9230 30405 9270
rect 30445 9230 30460 9270
rect 30390 8935 30460 9230
rect 30390 8900 30405 8935
rect 30445 8900 30460 8935
rect 30390 8640 30460 8900
rect 30390 8600 30405 8640
rect 30445 8600 30460 8640
rect 30390 8585 30460 8600
rect 31590 9270 31660 9285
rect 31590 9230 31605 9270
rect 31645 9230 31660 9270
rect 31590 8935 31660 9230
rect 32070 9270 32140 9285
rect 32070 9230 32085 9270
rect 32125 9230 32140 9270
rect 31590 8900 31605 8935
rect 31645 8900 31660 8935
rect 31590 8640 31660 8900
rect 31820 8670 31905 9200
rect 32070 8935 32140 9230
rect 32070 8900 32085 8935
rect 32125 8900 32140 8935
rect 31590 8600 31605 8640
rect 31645 8600 31660 8640
rect 31590 8585 31660 8600
rect 32070 8640 32140 8900
rect 32070 8600 32085 8640
rect 32125 8600 32140 8640
rect 32070 8585 32140 8600
rect 33270 9270 33340 9285
rect 33270 9230 33285 9270
rect 33325 9230 33340 9270
rect 33270 8935 33340 9230
rect 33270 8900 33285 8935
rect 33325 8900 33340 8935
rect 33270 8640 33340 8900
rect 33270 8600 33285 8640
rect 33325 8600 33340 8640
rect 33270 8585 33340 8600
rect 34325 8415 34400 9500
rect 35345 9270 35415 9285
rect 35345 9230 35360 9270
rect 35400 9230 35415 9270
rect 35345 8935 35415 9230
rect 35345 8900 35360 8935
rect 35400 8900 35415 8935
rect 35345 8640 35415 8900
rect 35345 8600 35360 8640
rect 35400 8600 35415 8640
rect 35345 8585 35415 8600
rect 36545 9270 36615 9285
rect 36545 9230 36560 9270
rect 36600 9230 36615 9270
rect 36545 8935 36615 9230
rect 37025 9270 37095 9285
rect 37025 9230 37040 9270
rect 37080 9230 37095 9270
rect 36545 8900 36560 8935
rect 36600 8900 36615 8935
rect 36545 8640 36615 8900
rect 36775 8670 36860 9200
rect 37025 8935 37095 9230
rect 37025 8900 37040 8935
rect 37080 8900 37095 8935
rect 36545 8600 36560 8640
rect 36600 8600 36615 8640
rect 36545 8585 36615 8600
rect 37025 8640 37095 8900
rect 37025 8600 37040 8640
rect 37080 8600 37095 8640
rect 37025 8585 37095 8600
rect 38225 9270 38295 9285
rect 38225 9230 38240 9270
rect 38280 9230 38295 9270
rect 38225 8935 38295 9230
rect 38225 8900 38240 8935
rect 38280 8900 38295 8935
rect 38225 8640 38295 8900
rect 38225 8600 38240 8640
rect 38280 8600 38295 8640
rect 38225 8585 38295 8600
rect 39280 8415 39355 9500
rect 40300 9270 40370 9285
rect 40300 9230 40315 9270
rect 40355 9230 40370 9270
rect 40300 8935 40370 9230
rect 40300 8900 40315 8935
rect 40355 8900 40370 8935
rect 40300 8640 40370 8900
rect 40300 8600 40315 8640
rect 40355 8600 40370 8640
rect 40300 8585 40370 8600
rect 41500 9270 41570 9285
rect 41500 9230 41515 9270
rect 41555 9230 41570 9270
rect 41500 8935 41570 9230
rect 41980 9270 42050 9285
rect 41980 9230 41995 9270
rect 42035 9230 42050 9270
rect 41500 8900 41515 8935
rect 41555 8900 41570 8935
rect 41500 8640 41570 8900
rect 41730 8670 41815 9200
rect 41980 8935 42050 9230
rect 41980 8900 41995 8935
rect 42035 8900 42050 8935
rect 41500 8600 41515 8640
rect 41555 8600 41570 8640
rect 41500 8585 41570 8600
rect 41980 8640 42050 8900
rect 41980 8600 41995 8640
rect 42035 8600 42050 8640
rect 41980 8585 42050 8600
rect 43180 9270 43250 9285
rect 43180 9230 43195 9270
rect 43235 9230 43250 9270
rect 43180 8935 43250 9230
rect 43180 8900 43195 8935
rect 43235 8900 43250 8935
rect 43180 8640 43250 8900
rect 43180 8600 43195 8640
rect 43235 8600 43250 8640
rect 43180 8585 43250 8600
rect 44235 8415 44310 9500
rect 45255 9270 45325 9285
rect 45255 9230 45270 9270
rect 45310 9230 45325 9270
rect 45255 8935 45325 9230
rect 45255 8900 45270 8935
rect 45310 8900 45325 8935
rect 45255 8640 45325 8900
rect 45255 8600 45270 8640
rect 45310 8600 45325 8640
rect 45255 8585 45325 8600
rect 46455 9270 46525 9285
rect 46455 9230 46470 9270
rect 46510 9230 46525 9270
rect 46455 8935 46525 9230
rect 46935 9270 47005 9285
rect 46935 9230 46950 9270
rect 46990 9230 47005 9270
rect 46455 8900 46470 8935
rect 46510 8900 46525 8935
rect 46455 8640 46525 8900
rect 46685 8670 46770 9200
rect 46935 8935 47005 9230
rect 46935 8900 46950 8935
rect 46990 8900 47005 8935
rect 46455 8600 46470 8640
rect 46510 8600 46525 8640
rect 46455 8585 46525 8600
rect 46935 8640 47005 8900
rect 46935 8600 46950 8640
rect 46990 8600 47005 8640
rect 46935 8585 47005 8600
rect 48135 9270 48205 9285
rect 48135 9230 48150 9270
rect 48190 9230 48205 9270
rect 48135 8935 48205 9230
rect 48135 8900 48150 8935
rect 48190 8900 48205 8935
rect 48135 8640 48205 8900
rect 48135 8600 48150 8640
rect 48190 8600 48205 8640
rect 48135 8585 48205 8600
rect 49190 8415 49265 9500
rect 50210 9270 50280 9285
rect 50210 9230 50225 9270
rect 50265 9230 50280 9270
rect 50210 8935 50280 9230
rect 50210 8900 50225 8935
rect 50265 8900 50280 8935
rect 50210 8640 50280 8900
rect 50210 8600 50225 8640
rect 50265 8600 50280 8640
rect 50210 8585 50280 8600
rect 51410 9270 51480 9285
rect 51410 9230 51425 9270
rect 51465 9230 51480 9270
rect 51410 8935 51480 9230
rect 51890 9270 51960 9285
rect 51890 9230 51905 9270
rect 51945 9230 51960 9270
rect 51410 8900 51425 8935
rect 51465 8900 51480 8935
rect 51410 8640 51480 8900
rect 51640 8670 51725 9200
rect 51890 8935 51960 9230
rect 51890 8900 51905 8935
rect 51945 8900 51960 8935
rect 51410 8600 51425 8640
rect 51465 8600 51480 8640
rect 51410 8585 51480 8600
rect 51890 8640 51960 8900
rect 51890 8600 51905 8640
rect 51945 8600 51960 8640
rect 51890 8585 51960 8600
rect 53090 9270 53160 9285
rect 53090 9230 53105 9270
rect 53145 9230 53160 9270
rect 53090 8935 53160 9230
rect 53090 8900 53105 8935
rect 53145 8900 53160 8935
rect 53090 8640 53160 8900
rect 53090 8600 53105 8640
rect 53145 8600 53160 8640
rect 53090 8585 53160 8600
rect 54145 8415 54220 9500
rect 55165 9270 55235 9285
rect 55165 9230 55180 9270
rect 55220 9230 55235 9270
rect 55165 8935 55235 9230
rect 55165 8900 55180 8935
rect 55220 8900 55235 8935
rect 55165 8640 55235 8900
rect 55165 8600 55180 8640
rect 55220 8600 55235 8640
rect 55165 8585 55235 8600
rect 56365 9270 56435 9285
rect 56365 9230 56380 9270
rect 56420 9230 56435 9270
rect 56365 8935 56435 9230
rect 56845 9270 56915 9285
rect 56845 9230 56860 9270
rect 56900 9230 56915 9270
rect 56365 8900 56380 8935
rect 56420 8900 56435 8935
rect 56365 8640 56435 8900
rect 56595 8670 56680 9200
rect 56845 8935 56915 9230
rect 56845 8900 56860 8935
rect 56900 8900 56915 8935
rect 56365 8600 56380 8640
rect 56420 8600 56435 8640
rect 56365 8585 56435 8600
rect 56845 8640 56915 8900
rect 56845 8600 56860 8640
rect 56900 8600 56915 8640
rect 56845 8585 56915 8600
rect 58045 9270 58115 9285
rect 58045 9230 58060 9270
rect 58100 9230 58115 9270
rect 58045 8935 58115 9230
rect 58045 8900 58060 8935
rect 58100 8900 58115 8935
rect 58045 8640 58115 8900
rect 58045 8600 58060 8640
rect 58100 8600 58115 8640
rect 58045 8585 58115 8600
rect 59100 8415 59175 9500
rect 60120 9270 60190 9285
rect 60120 9230 60135 9270
rect 60175 9230 60190 9270
rect 60120 8935 60190 9230
rect 60120 8900 60135 8935
rect 60175 8900 60190 8935
rect 60120 8640 60190 8900
rect 60120 8600 60135 8640
rect 60175 8600 60190 8640
rect 60120 8585 60190 8600
rect 61320 9270 61390 9285
rect 61320 9230 61335 9270
rect 61375 9230 61390 9270
rect 61320 8935 61390 9230
rect 61800 9270 61870 9285
rect 61800 9230 61815 9270
rect 61855 9230 61870 9270
rect 61320 8900 61335 8935
rect 61375 8900 61390 8935
rect 61320 8640 61390 8900
rect 61550 8670 61635 9200
rect 61800 8935 61870 9230
rect 61800 8900 61815 8935
rect 61855 8900 61870 8935
rect 61320 8600 61335 8640
rect 61375 8600 61390 8640
rect 61320 8585 61390 8600
rect 61800 8640 61870 8900
rect 61800 8600 61815 8640
rect 61855 8600 61870 8640
rect 61800 8585 61870 8600
rect 63000 9270 63070 9285
rect 63000 9230 63015 9270
rect 63055 9230 63070 9270
rect 63000 8935 63070 9230
rect 63000 8900 63015 8935
rect 63055 8900 63070 8935
rect 63000 8640 63070 8900
rect 63000 8600 63015 8640
rect 63055 8600 63070 8640
rect 63000 8585 63070 8600
rect 64055 8415 64130 9500
rect 65075 9270 65145 9285
rect 65075 9230 65090 9270
rect 65130 9230 65145 9270
rect 65075 8935 65145 9230
rect 65075 8900 65090 8935
rect 65130 8900 65145 8935
rect 65075 8640 65145 8900
rect 65075 8600 65090 8640
rect 65130 8600 65145 8640
rect 65075 8585 65145 8600
rect 66275 9270 66345 9285
rect 66275 9230 66290 9270
rect 66330 9230 66345 9270
rect 66275 8935 66345 9230
rect 66755 9270 66825 9285
rect 66755 9230 66770 9270
rect 66810 9230 66825 9270
rect 66275 8900 66290 8935
rect 66330 8900 66345 8935
rect 66275 8640 66345 8900
rect 66505 8670 66590 9200
rect 66755 8935 66825 9230
rect 66755 8900 66770 8935
rect 66810 8900 66825 8935
rect 66275 8600 66290 8640
rect 66330 8600 66345 8640
rect 66275 8585 66345 8600
rect 66755 8640 66825 8900
rect 66755 8600 66770 8640
rect 66810 8600 66825 8640
rect 66755 8585 66825 8600
rect 67955 9270 68025 9285
rect 67955 9230 67970 9270
rect 68010 9230 68025 9270
rect 67955 8935 68025 9230
rect 67955 8900 67970 8935
rect 68010 8900 68025 8935
rect 67955 8640 68025 8900
rect 67955 8600 67970 8640
rect 68010 8600 68025 8640
rect 67955 8585 68025 8600
rect 69010 8415 69085 9500
rect 70030 9270 70100 9285
rect 70030 9230 70045 9270
rect 70085 9230 70100 9270
rect 70030 8935 70100 9230
rect 70030 8900 70045 8935
rect 70085 8900 70100 8935
rect 70030 8640 70100 8900
rect 70030 8600 70045 8640
rect 70085 8600 70100 8640
rect 70030 8585 70100 8600
rect 71230 9270 71300 9285
rect 71230 9230 71245 9270
rect 71285 9230 71300 9270
rect 71230 8935 71300 9230
rect 71710 9270 71780 9285
rect 71710 9230 71725 9270
rect 71765 9230 71780 9270
rect 71230 8900 71245 8935
rect 71285 8900 71300 8935
rect 71230 8640 71300 8900
rect 71460 8670 71545 9200
rect 71710 8935 71780 9230
rect 71710 8900 71725 8935
rect 71765 8900 71780 8935
rect 71230 8600 71245 8640
rect 71285 8600 71300 8640
rect 71230 8585 71300 8600
rect 71710 8640 71780 8900
rect 71710 8600 71725 8640
rect 71765 8600 71780 8640
rect 71710 8585 71780 8600
rect 72910 9270 72980 9285
rect 72910 9230 72925 9270
rect 72965 9230 72980 9270
rect 72910 8935 72980 9230
rect 72910 8900 72925 8935
rect 72965 8900 72980 8935
rect 72910 8640 72980 8900
rect 72910 8600 72925 8640
rect 72965 8600 72980 8640
rect 72910 8585 72980 8600
rect 73965 8415 74040 9500
rect 74985 9270 75055 9285
rect 74985 9230 75000 9270
rect 75040 9230 75055 9270
rect 74985 8935 75055 9230
rect 74985 8900 75000 8935
rect 75040 8900 75055 8935
rect 74985 8640 75055 8900
rect 74985 8600 75000 8640
rect 75040 8600 75055 8640
rect 74985 8585 75055 8600
rect 76185 9270 76255 9285
rect 76185 9230 76200 9270
rect 76240 9230 76255 9270
rect 76185 8935 76255 9230
rect 76665 9270 76735 9285
rect 76665 9230 76680 9270
rect 76720 9230 76735 9270
rect 76185 8900 76200 8935
rect 76240 8900 76255 8935
rect 76185 8640 76255 8900
rect 76415 8670 76500 9200
rect 76665 8935 76735 9230
rect 76665 8900 76680 8935
rect 76720 8900 76735 8935
rect 76185 8600 76200 8640
rect 76240 8600 76255 8640
rect 76185 8585 76255 8600
rect 76665 8640 76735 8900
rect 76665 8600 76680 8640
rect 76720 8600 76735 8640
rect 76665 8585 76735 8600
rect 77865 9270 77935 9285
rect 77865 9230 77880 9270
rect 77920 9230 77935 9270
rect 77865 8935 77935 9230
rect 77865 8900 77880 8935
rect 77920 8900 77935 8935
rect 77865 8640 77935 8900
rect 77865 8600 77880 8640
rect 77920 8600 77935 8640
rect 77865 8585 77935 8600
rect 3735 8345 5485 8415
rect 8690 8400 10440 8415
rect 8690 8360 8705 8400
rect 8745 8360 10385 8400
rect 10425 8360 10440 8400
rect 8690 8345 10440 8360
rect 13645 8400 15395 8415
rect 13645 8360 13660 8400
rect 13700 8360 15340 8400
rect 15380 8360 15395 8400
rect 13645 8345 15395 8360
rect 18600 8400 20350 8415
rect 18600 8360 18615 8400
rect 18655 8360 20295 8400
rect 20335 8360 20350 8400
rect 18600 8345 20350 8360
rect 23555 8400 25305 8415
rect 23555 8360 23570 8400
rect 23610 8360 25250 8400
rect 25290 8360 25305 8400
rect 23555 8345 25305 8360
rect 28510 8400 30260 8415
rect 28510 8360 28525 8400
rect 28565 8360 30205 8400
rect 30245 8360 30260 8400
rect 28510 8345 30260 8360
rect 33465 8400 35215 8415
rect 33465 8360 33480 8400
rect 33520 8360 35160 8400
rect 35200 8360 35215 8400
rect 33465 8345 35215 8360
rect 38420 8400 40170 8415
rect 38420 8360 38435 8400
rect 38475 8360 40115 8400
rect 40155 8360 40170 8400
rect 38420 8345 40170 8360
rect 43375 8400 45125 8415
rect 43375 8360 43390 8400
rect 43430 8360 45070 8400
rect 45110 8360 45125 8400
rect 43375 8345 45125 8360
rect 48330 8400 50080 8415
rect 48330 8360 48345 8400
rect 48385 8360 50025 8400
rect 50065 8360 50080 8400
rect 48330 8345 50080 8360
rect 53285 8400 55035 8415
rect 53285 8360 53300 8400
rect 53340 8360 54980 8400
rect 55020 8360 55035 8400
rect 53285 8345 55035 8360
rect 58240 8400 59990 8415
rect 58240 8360 58255 8400
rect 58295 8360 59935 8400
rect 59975 8360 59990 8400
rect 58240 8345 59990 8360
rect 63195 8400 64945 8415
rect 63195 8360 63210 8400
rect 63250 8360 64890 8400
rect 64930 8360 64945 8400
rect 63195 8345 64945 8360
rect 68150 8400 69900 8415
rect 68150 8360 68165 8400
rect 68205 8360 69845 8400
rect 69885 8360 69900 8400
rect 68150 8345 69900 8360
rect 73105 8400 74855 8415
rect 73105 8360 73120 8400
rect 73160 8360 74800 8400
rect 74840 8360 74855 8400
rect 73105 8345 74855 8360
rect 4595 6495 4670 8345
rect 9550 6495 9625 8345
rect 14505 6495 14580 8345
rect 19460 6495 19535 8345
rect 24415 6495 24490 8345
rect 29370 6495 29445 8345
rect 34325 6495 34400 8345
rect 39280 6495 39355 8345
rect 44235 6495 44310 8345
rect 49190 6495 49265 8345
rect 54145 6495 54220 8345
rect 59100 6495 59175 8345
rect 64055 6495 64130 8345
rect 69010 6495 69085 8345
rect 73965 6495 74040 8345
rect 3735 6425 5485 6495
rect 8690 6480 10440 6495
rect 8690 6440 8705 6480
rect 8745 6440 10385 6480
rect 10425 6440 10440 6480
rect 8690 6425 10440 6440
rect 13645 6480 15395 6495
rect 13645 6440 13660 6480
rect 13700 6440 15340 6480
rect 15380 6440 15395 6480
rect 13645 6425 15395 6440
rect 18600 6480 20350 6495
rect 18600 6440 18615 6480
rect 18655 6440 20295 6480
rect 20335 6440 20350 6480
rect 18600 6425 20350 6440
rect 23555 6480 25305 6495
rect 23555 6440 23570 6480
rect 23610 6440 25250 6480
rect 25290 6440 25305 6480
rect 23555 6425 25305 6440
rect 28510 6480 30260 6495
rect 28510 6440 28525 6480
rect 28565 6440 30205 6480
rect 30245 6440 30260 6480
rect 28510 6425 30260 6440
rect 33465 6480 35215 6495
rect 33465 6440 33480 6480
rect 33520 6440 35160 6480
rect 35200 6440 35215 6480
rect 33465 6425 35215 6440
rect 38420 6480 40170 6495
rect 38420 6440 38435 6480
rect 38475 6440 40115 6480
rect 40155 6440 40170 6480
rect 38420 6425 40170 6440
rect 43375 6480 45125 6495
rect 43375 6440 43390 6480
rect 43430 6440 45070 6480
rect 45110 6440 45125 6480
rect 43375 6425 45125 6440
rect 48330 6480 50080 6495
rect 48330 6440 48345 6480
rect 48385 6440 50025 6480
rect 50065 6440 50080 6480
rect 48330 6425 50080 6440
rect 53285 6480 55035 6495
rect 53285 6440 53300 6480
rect 53340 6440 54980 6480
rect 55020 6440 55035 6480
rect 53285 6425 55035 6440
rect 58240 6480 59990 6495
rect 58240 6440 58255 6480
rect 58295 6440 59935 6480
rect 59975 6440 59990 6480
rect 58240 6425 59990 6440
rect 63195 6480 64945 6495
rect 63195 6440 63210 6480
rect 63250 6440 64890 6480
rect 64930 6440 64945 6480
rect 63195 6425 64945 6440
rect 68150 6480 69900 6495
rect 68150 6440 68165 6480
rect 68205 6440 69845 6480
rect 69885 6440 69900 6480
rect 68150 6425 69900 6440
rect 73105 6480 74855 6495
rect 73105 6440 73120 6480
rect 73160 6440 74800 6480
rect 74840 6440 74855 6480
rect 73105 6425 74855 6440
rect 660 5885 730 6210
rect 660 5850 675 5885
rect 715 5850 730 5885
rect 660 5510 730 5850
rect 1860 5885 1930 6210
rect 1860 5850 1875 5885
rect 1915 5850 1930 5885
rect 1860 5510 1930 5850
rect 2090 5595 2175 6125
rect 2340 5885 2410 6210
rect 2340 5850 2355 5885
rect 2395 5850 2410 5885
rect 2340 5510 2410 5850
rect 3540 5885 3610 6210
rect 3540 5850 3555 5885
rect 3595 5850 3610 5885
rect 3540 5510 3610 5850
rect 4595 5340 4670 6425
rect 5615 6195 5685 6210
rect 5615 6155 5630 6195
rect 5670 6155 5685 6195
rect 5615 5885 5685 6155
rect 5615 5850 5630 5885
rect 5670 5850 5685 5885
rect 5615 5565 5685 5850
rect 5615 5525 5630 5565
rect 5670 5525 5685 5565
rect 5615 5510 5685 5525
rect 6815 6195 6885 6210
rect 6815 6155 6830 6195
rect 6870 6155 6885 6195
rect 6815 5885 6885 6155
rect 7295 6195 7365 6210
rect 7295 6155 7310 6195
rect 7350 6155 7365 6195
rect 6815 5850 6830 5885
rect 6870 5850 6885 5885
rect 6815 5565 6885 5850
rect 7045 5595 7130 6125
rect 7295 5885 7365 6155
rect 7295 5850 7310 5885
rect 7350 5850 7365 5885
rect 6815 5525 6830 5565
rect 6870 5525 6885 5565
rect 6815 5510 6885 5525
rect 7295 5565 7365 5850
rect 7295 5525 7310 5565
rect 7350 5525 7365 5565
rect 7295 5510 7365 5525
rect 8495 6195 8565 6210
rect 8495 6155 8510 6195
rect 8550 6155 8565 6195
rect 8495 5885 8565 6155
rect 8495 5850 8510 5885
rect 8550 5850 8565 5885
rect 8495 5565 8565 5850
rect 8495 5525 8510 5565
rect 8550 5525 8565 5565
rect 8495 5510 8565 5525
rect 9550 5340 9625 6425
rect 10570 6195 10640 6210
rect 10570 6155 10585 6195
rect 10625 6155 10640 6195
rect 10570 5885 10640 6155
rect 10570 5850 10585 5885
rect 10625 5850 10640 5885
rect 10570 5565 10640 5850
rect 10570 5525 10585 5565
rect 10625 5525 10640 5565
rect 10570 5510 10640 5525
rect 11770 6195 11840 6210
rect 11770 6155 11785 6195
rect 11825 6155 11840 6195
rect 11770 5885 11840 6155
rect 12250 6195 12320 6210
rect 12250 6155 12265 6195
rect 12305 6155 12320 6195
rect 11770 5850 11785 5885
rect 11825 5850 11840 5885
rect 11770 5565 11840 5850
rect 12000 5595 12085 6125
rect 12250 5885 12320 6155
rect 12250 5850 12265 5885
rect 12305 5850 12320 5885
rect 11770 5525 11785 5565
rect 11825 5525 11840 5565
rect 11770 5510 11840 5525
rect 12250 5565 12320 5850
rect 12250 5525 12265 5565
rect 12305 5525 12320 5565
rect 12250 5510 12320 5525
rect 13450 6195 13520 6210
rect 13450 6155 13465 6195
rect 13505 6155 13520 6195
rect 13450 5885 13520 6155
rect 13450 5850 13465 5885
rect 13505 5850 13520 5885
rect 13450 5565 13520 5850
rect 13450 5525 13465 5565
rect 13505 5525 13520 5565
rect 13450 5510 13520 5525
rect 14505 5340 14580 6425
rect 15525 6195 15595 6210
rect 15525 6155 15540 6195
rect 15580 6155 15595 6195
rect 15525 5885 15595 6155
rect 15525 5850 15540 5885
rect 15580 5850 15595 5885
rect 15525 5565 15595 5850
rect 15525 5525 15540 5565
rect 15580 5525 15595 5565
rect 15525 5510 15595 5525
rect 16725 6195 16795 6210
rect 16725 6155 16740 6195
rect 16780 6155 16795 6195
rect 16725 5885 16795 6155
rect 17205 6195 17275 6210
rect 17205 6155 17220 6195
rect 17260 6155 17275 6195
rect 16725 5850 16740 5885
rect 16780 5850 16795 5885
rect 16725 5565 16795 5850
rect 16955 5595 17040 6125
rect 17205 5885 17275 6155
rect 17205 5850 17220 5885
rect 17260 5850 17275 5885
rect 16725 5525 16740 5565
rect 16780 5525 16795 5565
rect 16725 5510 16795 5525
rect 17205 5565 17275 5850
rect 17205 5525 17220 5565
rect 17260 5525 17275 5565
rect 17205 5510 17275 5525
rect 18405 6195 18475 6210
rect 18405 6155 18420 6195
rect 18460 6155 18475 6195
rect 18405 5885 18475 6155
rect 18405 5850 18420 5885
rect 18460 5850 18475 5885
rect 18405 5565 18475 5850
rect 18405 5525 18420 5565
rect 18460 5525 18475 5565
rect 18405 5510 18475 5525
rect 19460 5340 19535 6425
rect 20480 6195 20550 6210
rect 20480 6155 20495 6195
rect 20535 6155 20550 6195
rect 20480 5885 20550 6155
rect 20480 5850 20495 5885
rect 20535 5850 20550 5885
rect 20480 5565 20550 5850
rect 20480 5525 20495 5565
rect 20535 5525 20550 5565
rect 20480 5510 20550 5525
rect 21680 6195 21750 6210
rect 21680 6155 21695 6195
rect 21735 6155 21750 6195
rect 21680 5885 21750 6155
rect 22160 6195 22230 6210
rect 22160 6155 22175 6195
rect 22215 6155 22230 6195
rect 21680 5850 21695 5885
rect 21735 5850 21750 5885
rect 21680 5565 21750 5850
rect 21910 5595 21995 6125
rect 22160 5885 22230 6155
rect 22160 5850 22175 5885
rect 22215 5850 22230 5885
rect 21680 5525 21695 5565
rect 21735 5525 21750 5565
rect 21680 5510 21750 5525
rect 22160 5565 22230 5850
rect 22160 5525 22175 5565
rect 22215 5525 22230 5565
rect 22160 5510 22230 5525
rect 23360 6195 23430 6210
rect 23360 6155 23375 6195
rect 23415 6155 23430 6195
rect 23360 5885 23430 6155
rect 23360 5850 23375 5885
rect 23415 5850 23430 5885
rect 23360 5565 23430 5850
rect 23360 5525 23375 5565
rect 23415 5525 23430 5565
rect 23360 5510 23430 5525
rect 24415 5340 24490 6425
rect 25435 6195 25505 6210
rect 25435 6155 25450 6195
rect 25490 6155 25505 6195
rect 25435 5885 25505 6155
rect 25435 5850 25450 5885
rect 25490 5850 25505 5885
rect 25435 5565 25505 5850
rect 25435 5525 25450 5565
rect 25490 5525 25505 5565
rect 25435 5510 25505 5525
rect 26635 6195 26705 6210
rect 26635 6155 26650 6195
rect 26690 6155 26705 6195
rect 26635 5885 26705 6155
rect 27115 6195 27185 6210
rect 27115 6155 27130 6195
rect 27170 6155 27185 6195
rect 26635 5850 26650 5885
rect 26690 5850 26705 5885
rect 26635 5565 26705 5850
rect 26865 5595 26950 6125
rect 27115 5885 27185 6155
rect 27115 5850 27130 5885
rect 27170 5850 27185 5885
rect 26635 5525 26650 5565
rect 26690 5525 26705 5565
rect 26635 5510 26705 5525
rect 27115 5565 27185 5850
rect 27115 5525 27130 5565
rect 27170 5525 27185 5565
rect 27115 5510 27185 5525
rect 28315 6195 28385 6210
rect 28315 6155 28330 6195
rect 28370 6155 28385 6195
rect 28315 5885 28385 6155
rect 28315 5850 28330 5885
rect 28370 5850 28385 5885
rect 28315 5565 28385 5850
rect 28315 5525 28330 5565
rect 28370 5525 28385 5565
rect 28315 5510 28385 5525
rect 29370 5340 29445 6425
rect 30390 6195 30460 6210
rect 30390 6155 30405 6195
rect 30445 6155 30460 6195
rect 30390 5885 30460 6155
rect 30390 5850 30405 5885
rect 30445 5850 30460 5885
rect 30390 5565 30460 5850
rect 30390 5525 30405 5565
rect 30445 5525 30460 5565
rect 30390 5510 30460 5525
rect 31590 6195 31660 6210
rect 31590 6155 31605 6195
rect 31645 6155 31660 6195
rect 31590 5885 31660 6155
rect 32070 6195 32140 6210
rect 32070 6155 32085 6195
rect 32125 6155 32140 6195
rect 31590 5850 31605 5885
rect 31645 5850 31660 5885
rect 31590 5565 31660 5850
rect 31820 5595 31905 6125
rect 32070 5885 32140 6155
rect 32070 5850 32085 5885
rect 32125 5850 32140 5885
rect 31590 5525 31605 5565
rect 31645 5525 31660 5565
rect 31590 5510 31660 5525
rect 32070 5565 32140 5850
rect 32070 5525 32085 5565
rect 32125 5525 32140 5565
rect 32070 5510 32140 5525
rect 33270 6195 33340 6210
rect 33270 6155 33285 6195
rect 33325 6155 33340 6195
rect 33270 5885 33340 6155
rect 33270 5850 33285 5885
rect 33325 5850 33340 5885
rect 33270 5565 33340 5850
rect 33270 5525 33285 5565
rect 33325 5525 33340 5565
rect 33270 5510 33340 5525
rect 34325 5340 34400 6425
rect 35345 6195 35415 6210
rect 35345 6155 35360 6195
rect 35400 6155 35415 6195
rect 35345 5885 35415 6155
rect 35345 5850 35360 5885
rect 35400 5850 35415 5885
rect 35345 5565 35415 5850
rect 35345 5525 35360 5565
rect 35400 5525 35415 5565
rect 35345 5510 35415 5525
rect 36545 6195 36615 6210
rect 36545 6155 36560 6195
rect 36600 6155 36615 6195
rect 36545 5885 36615 6155
rect 37025 6195 37095 6210
rect 37025 6155 37040 6195
rect 37080 6155 37095 6195
rect 36545 5850 36560 5885
rect 36600 5850 36615 5885
rect 36545 5565 36615 5850
rect 36775 5595 36860 6125
rect 37025 5885 37095 6155
rect 37025 5850 37040 5885
rect 37080 5850 37095 5885
rect 36545 5525 36560 5565
rect 36600 5525 36615 5565
rect 36545 5510 36615 5525
rect 37025 5565 37095 5850
rect 37025 5525 37040 5565
rect 37080 5525 37095 5565
rect 37025 5510 37095 5525
rect 38225 6195 38295 6210
rect 38225 6155 38240 6195
rect 38280 6155 38295 6195
rect 38225 5885 38295 6155
rect 38225 5850 38240 5885
rect 38280 5850 38295 5885
rect 38225 5565 38295 5850
rect 38225 5525 38240 5565
rect 38280 5525 38295 5565
rect 38225 5510 38295 5525
rect 39280 5340 39355 6425
rect 40300 6195 40370 6210
rect 40300 6155 40315 6195
rect 40355 6155 40370 6195
rect 40300 5885 40370 6155
rect 40300 5850 40315 5885
rect 40355 5850 40370 5885
rect 40300 5565 40370 5850
rect 40300 5525 40315 5565
rect 40355 5525 40370 5565
rect 40300 5510 40370 5525
rect 41500 6195 41570 6210
rect 41500 6155 41515 6195
rect 41555 6155 41570 6195
rect 41500 5885 41570 6155
rect 41980 6195 42050 6210
rect 41980 6155 41995 6195
rect 42035 6155 42050 6195
rect 41500 5850 41515 5885
rect 41555 5850 41570 5885
rect 41500 5565 41570 5850
rect 41730 5595 41815 6125
rect 41980 5885 42050 6155
rect 41980 5850 41995 5885
rect 42035 5850 42050 5885
rect 41500 5525 41515 5565
rect 41555 5525 41570 5565
rect 41500 5510 41570 5525
rect 41980 5565 42050 5850
rect 41980 5525 41995 5565
rect 42035 5525 42050 5565
rect 41980 5510 42050 5525
rect 43180 6195 43250 6210
rect 43180 6155 43195 6195
rect 43235 6155 43250 6195
rect 43180 5885 43250 6155
rect 43180 5850 43195 5885
rect 43235 5850 43250 5885
rect 43180 5565 43250 5850
rect 43180 5525 43195 5565
rect 43235 5525 43250 5565
rect 43180 5510 43250 5525
rect 44235 5340 44310 6425
rect 45255 6195 45325 6210
rect 45255 6155 45270 6195
rect 45310 6155 45325 6195
rect 45255 5885 45325 6155
rect 45255 5850 45270 5885
rect 45310 5850 45325 5885
rect 45255 5565 45325 5850
rect 45255 5525 45270 5565
rect 45310 5525 45325 5565
rect 45255 5510 45325 5525
rect 46455 6195 46525 6210
rect 46455 6155 46470 6195
rect 46510 6155 46525 6195
rect 46455 5885 46525 6155
rect 46935 6195 47005 6210
rect 46935 6155 46950 6195
rect 46990 6155 47005 6195
rect 46455 5850 46470 5885
rect 46510 5850 46525 5885
rect 46455 5565 46525 5850
rect 46685 5595 46770 6125
rect 46935 5885 47005 6155
rect 46935 5850 46950 5885
rect 46990 5850 47005 5885
rect 46455 5525 46470 5565
rect 46510 5525 46525 5565
rect 46455 5510 46525 5525
rect 46935 5565 47005 5850
rect 46935 5525 46950 5565
rect 46990 5525 47005 5565
rect 46935 5510 47005 5525
rect 48135 6195 48205 6210
rect 48135 6155 48150 6195
rect 48190 6155 48205 6195
rect 48135 5885 48205 6155
rect 48135 5850 48150 5885
rect 48190 5850 48205 5885
rect 48135 5565 48205 5850
rect 48135 5525 48150 5565
rect 48190 5525 48205 5565
rect 48135 5510 48205 5525
rect 49190 5340 49265 6425
rect 50210 6195 50280 6210
rect 50210 6155 50225 6195
rect 50265 6155 50280 6195
rect 50210 5885 50280 6155
rect 50210 5850 50225 5885
rect 50265 5850 50280 5885
rect 50210 5565 50280 5850
rect 50210 5525 50225 5565
rect 50265 5525 50280 5565
rect 50210 5510 50280 5525
rect 51410 6195 51480 6210
rect 51410 6155 51425 6195
rect 51465 6155 51480 6195
rect 51410 5885 51480 6155
rect 51890 6195 51960 6210
rect 51890 6155 51905 6195
rect 51945 6155 51960 6195
rect 51410 5850 51425 5885
rect 51465 5850 51480 5885
rect 51410 5565 51480 5850
rect 51640 5595 51725 6125
rect 51890 5885 51960 6155
rect 51890 5850 51905 5885
rect 51945 5850 51960 5885
rect 51410 5525 51425 5565
rect 51465 5525 51480 5565
rect 51410 5510 51480 5525
rect 51890 5565 51960 5850
rect 51890 5525 51905 5565
rect 51945 5525 51960 5565
rect 51890 5510 51960 5525
rect 53090 6195 53160 6210
rect 53090 6155 53105 6195
rect 53145 6155 53160 6195
rect 53090 5885 53160 6155
rect 53090 5850 53105 5885
rect 53145 5850 53160 5885
rect 53090 5565 53160 5850
rect 53090 5525 53105 5565
rect 53145 5525 53160 5565
rect 53090 5510 53160 5525
rect 54145 5340 54220 6425
rect 55165 6195 55235 6210
rect 55165 6155 55180 6195
rect 55220 6155 55235 6195
rect 55165 5885 55235 6155
rect 55165 5850 55180 5885
rect 55220 5850 55235 5885
rect 55165 5565 55235 5850
rect 55165 5525 55180 5565
rect 55220 5525 55235 5565
rect 55165 5510 55235 5525
rect 56365 6195 56435 6210
rect 56365 6155 56380 6195
rect 56420 6155 56435 6195
rect 56365 5885 56435 6155
rect 56845 6195 56915 6210
rect 56845 6155 56860 6195
rect 56900 6155 56915 6195
rect 56365 5850 56380 5885
rect 56420 5850 56435 5885
rect 56365 5565 56435 5850
rect 56595 5595 56680 6125
rect 56845 5885 56915 6155
rect 56845 5850 56860 5885
rect 56900 5850 56915 5885
rect 56365 5525 56380 5565
rect 56420 5525 56435 5565
rect 56365 5510 56435 5525
rect 56845 5565 56915 5850
rect 56845 5525 56860 5565
rect 56900 5525 56915 5565
rect 56845 5510 56915 5525
rect 58045 6195 58115 6210
rect 58045 6155 58060 6195
rect 58100 6155 58115 6195
rect 58045 5885 58115 6155
rect 58045 5850 58060 5885
rect 58100 5850 58115 5885
rect 58045 5565 58115 5850
rect 58045 5525 58060 5565
rect 58100 5525 58115 5565
rect 58045 5510 58115 5525
rect 59100 5340 59175 6425
rect 60120 6195 60190 6210
rect 60120 6155 60135 6195
rect 60175 6155 60190 6195
rect 60120 5885 60190 6155
rect 60120 5850 60135 5885
rect 60175 5850 60190 5885
rect 60120 5565 60190 5850
rect 60120 5525 60135 5565
rect 60175 5525 60190 5565
rect 60120 5510 60190 5525
rect 61320 6195 61390 6210
rect 61320 6155 61335 6195
rect 61375 6155 61390 6195
rect 61320 5885 61390 6155
rect 61800 6195 61870 6210
rect 61800 6155 61815 6195
rect 61855 6155 61870 6195
rect 61320 5850 61335 5885
rect 61375 5850 61390 5885
rect 61320 5565 61390 5850
rect 61550 5595 61635 6125
rect 61800 5885 61870 6155
rect 61800 5850 61815 5885
rect 61855 5850 61870 5885
rect 61320 5525 61335 5565
rect 61375 5525 61390 5565
rect 61320 5510 61390 5525
rect 61800 5565 61870 5850
rect 61800 5525 61815 5565
rect 61855 5525 61870 5565
rect 61800 5510 61870 5525
rect 63000 6195 63070 6210
rect 63000 6155 63015 6195
rect 63055 6155 63070 6195
rect 63000 5885 63070 6155
rect 63000 5850 63015 5885
rect 63055 5850 63070 5885
rect 63000 5565 63070 5850
rect 63000 5525 63015 5565
rect 63055 5525 63070 5565
rect 63000 5510 63070 5525
rect 64055 5340 64130 6425
rect 65075 6195 65145 6210
rect 65075 6155 65090 6195
rect 65130 6155 65145 6195
rect 65075 5885 65145 6155
rect 65075 5850 65090 5885
rect 65130 5850 65145 5885
rect 65075 5565 65145 5850
rect 65075 5525 65090 5565
rect 65130 5525 65145 5565
rect 65075 5510 65145 5525
rect 66275 6195 66345 6210
rect 66275 6155 66290 6195
rect 66330 6155 66345 6195
rect 66275 5885 66345 6155
rect 66755 6195 66825 6210
rect 66755 6155 66770 6195
rect 66810 6155 66825 6195
rect 66275 5850 66290 5885
rect 66330 5850 66345 5885
rect 66275 5565 66345 5850
rect 66505 5595 66590 6125
rect 66755 5885 66825 6155
rect 66755 5850 66770 5885
rect 66810 5850 66825 5885
rect 66275 5525 66290 5565
rect 66330 5525 66345 5565
rect 66275 5510 66345 5525
rect 66755 5565 66825 5850
rect 66755 5525 66770 5565
rect 66810 5525 66825 5565
rect 66755 5510 66825 5525
rect 67955 6195 68025 6210
rect 67955 6155 67970 6195
rect 68010 6155 68025 6195
rect 67955 5885 68025 6155
rect 67955 5850 67970 5885
rect 68010 5850 68025 5885
rect 67955 5565 68025 5850
rect 67955 5525 67970 5565
rect 68010 5525 68025 5565
rect 67955 5510 68025 5525
rect 69010 5340 69085 6425
rect 70030 6195 70100 6210
rect 70030 6155 70045 6195
rect 70085 6155 70100 6195
rect 70030 5885 70100 6155
rect 70030 5850 70045 5885
rect 70085 5850 70100 5885
rect 70030 5565 70100 5850
rect 70030 5525 70045 5565
rect 70085 5525 70100 5565
rect 70030 5510 70100 5525
rect 71230 6195 71300 6210
rect 71230 6155 71245 6195
rect 71285 6155 71300 6195
rect 71230 5885 71300 6155
rect 71710 6195 71780 6210
rect 71710 6155 71725 6195
rect 71765 6155 71780 6195
rect 71230 5850 71245 5885
rect 71285 5850 71300 5885
rect 71230 5565 71300 5850
rect 71460 5595 71545 6125
rect 71710 5885 71780 6155
rect 71710 5850 71725 5885
rect 71765 5850 71780 5885
rect 71230 5525 71245 5565
rect 71285 5525 71300 5565
rect 71230 5510 71300 5525
rect 71710 5565 71780 5850
rect 71710 5525 71725 5565
rect 71765 5525 71780 5565
rect 71710 5510 71780 5525
rect 72910 6195 72980 6210
rect 72910 6155 72925 6195
rect 72965 6155 72980 6195
rect 72910 5885 72980 6155
rect 72910 5850 72925 5885
rect 72965 5850 72980 5885
rect 72910 5565 72980 5850
rect 72910 5525 72925 5565
rect 72965 5525 72980 5565
rect 72910 5510 72980 5525
rect 73965 5340 74040 6425
rect 74985 6195 75055 6210
rect 74985 6155 75000 6195
rect 75040 6155 75055 6195
rect 74985 5885 75055 6155
rect 74985 5850 75000 5885
rect 75040 5850 75055 5885
rect 74985 5565 75055 5850
rect 74985 5525 75000 5565
rect 75040 5525 75055 5565
rect 74985 5510 75055 5525
rect 76185 6195 76255 6210
rect 76185 6155 76200 6195
rect 76240 6155 76255 6195
rect 76185 5885 76255 6155
rect 76665 6195 76735 6210
rect 76665 6155 76680 6195
rect 76720 6155 76735 6195
rect 76185 5850 76200 5885
rect 76240 5850 76255 5885
rect 76185 5565 76255 5850
rect 76415 5595 76500 6125
rect 76665 5885 76735 6155
rect 76665 5850 76680 5885
rect 76720 5850 76735 5885
rect 76185 5525 76200 5565
rect 76240 5525 76255 5565
rect 76185 5510 76255 5525
rect 76665 5565 76735 5850
rect 76665 5525 76680 5565
rect 76720 5525 76735 5565
rect 76665 5510 76735 5525
rect 77865 6195 77935 6210
rect 77865 6155 77880 6195
rect 77920 6155 77935 6195
rect 77865 5885 77935 6155
rect 77865 5850 77880 5885
rect 77920 5850 77935 5885
rect 77865 5565 77935 5850
rect 77865 5525 77880 5565
rect 77920 5525 77935 5565
rect 77865 5510 77935 5525
rect 3735 5270 5485 5340
rect 8690 5325 10440 5340
rect 8690 5285 8705 5325
rect 8745 5285 10385 5325
rect 10425 5285 10440 5325
rect 8690 5270 10440 5285
rect 13645 5325 15395 5340
rect 13645 5285 13660 5325
rect 13700 5285 15340 5325
rect 15380 5285 15395 5325
rect 13645 5270 15395 5285
rect 18600 5325 20350 5340
rect 18600 5285 18615 5325
rect 18655 5285 20295 5325
rect 20335 5285 20350 5325
rect 18600 5270 20350 5285
rect 23555 5325 25305 5340
rect 23555 5285 23570 5325
rect 23610 5285 25250 5325
rect 25290 5285 25305 5325
rect 23555 5270 25305 5285
rect 28510 5325 30260 5340
rect 28510 5285 28525 5325
rect 28565 5285 30205 5325
rect 30245 5285 30260 5325
rect 28510 5270 30260 5285
rect 33465 5325 35215 5340
rect 33465 5285 33480 5325
rect 33520 5285 35160 5325
rect 35200 5285 35215 5325
rect 33465 5270 35215 5285
rect 38420 5325 40170 5340
rect 38420 5285 38435 5325
rect 38475 5285 40115 5325
rect 40155 5285 40170 5325
rect 38420 5270 40170 5285
rect 43375 5325 45125 5340
rect 43375 5285 43390 5325
rect 43430 5285 45070 5325
rect 45110 5285 45125 5325
rect 43375 5270 45125 5285
rect 48330 5325 50080 5340
rect 48330 5285 48345 5325
rect 48385 5285 50025 5325
rect 50065 5285 50080 5325
rect 48330 5270 50080 5285
rect 53285 5325 55035 5340
rect 53285 5285 53300 5325
rect 53340 5285 54980 5325
rect 55020 5285 55035 5325
rect 53285 5270 55035 5285
rect 58240 5325 59990 5340
rect 58240 5285 58255 5325
rect 58295 5285 59935 5325
rect 59975 5285 59990 5325
rect 58240 5270 59990 5285
rect 63195 5325 64945 5340
rect 63195 5285 63210 5325
rect 63250 5285 64890 5325
rect 64930 5285 64945 5325
rect 63195 5270 64945 5285
rect 68150 5325 69900 5340
rect 68150 5285 68165 5325
rect 68205 5285 69845 5325
rect 69885 5285 69900 5325
rect 68150 5270 69900 5285
rect 73105 5325 74855 5340
rect 73105 5285 73120 5325
rect 73160 5285 74800 5325
rect 74840 5285 74855 5325
rect 73105 5270 74855 5285
rect 4595 3420 4670 5270
rect 9550 3420 9625 5270
rect 14505 3420 14580 5270
rect 19460 3420 19535 5270
rect 24415 3420 24490 5270
rect 29370 3420 29445 5270
rect 34325 3420 34400 5270
rect 39280 3420 39355 5270
rect 44235 3420 44310 5270
rect 49190 3420 49265 5270
rect 54145 3420 54220 5270
rect 59100 3420 59175 5270
rect 64055 3420 64130 5270
rect 69010 3420 69085 5270
rect 73965 3420 74040 5270
rect 3735 3350 5485 3420
rect 8690 3405 10440 3420
rect 8690 3365 8705 3405
rect 8745 3365 10385 3405
rect 10425 3365 10440 3405
rect 8690 3350 10440 3365
rect 13645 3405 15395 3420
rect 13645 3365 13660 3405
rect 13700 3365 15340 3405
rect 15380 3365 15395 3405
rect 13645 3350 15395 3365
rect 18600 3405 20350 3420
rect 18600 3365 18615 3405
rect 18655 3365 20295 3405
rect 20335 3365 20350 3405
rect 18600 3350 20350 3365
rect 23555 3405 25305 3420
rect 23555 3365 23570 3405
rect 23610 3365 25250 3405
rect 25290 3365 25305 3405
rect 23555 3350 25305 3365
rect 28510 3405 30260 3420
rect 28510 3365 28525 3405
rect 28565 3365 30205 3405
rect 30245 3365 30260 3405
rect 28510 3350 30260 3365
rect 33465 3405 35215 3420
rect 33465 3365 33480 3405
rect 33520 3365 35160 3405
rect 35200 3365 35215 3405
rect 33465 3350 35215 3365
rect 38420 3405 40170 3420
rect 38420 3365 38435 3405
rect 38475 3365 40115 3405
rect 40155 3365 40170 3405
rect 38420 3350 40170 3365
rect 43375 3405 45125 3420
rect 43375 3365 43390 3405
rect 43430 3365 45070 3405
rect 45110 3365 45125 3405
rect 43375 3350 45125 3365
rect 48330 3405 50080 3420
rect 48330 3365 48345 3405
rect 48385 3365 50025 3405
rect 50065 3365 50080 3405
rect 48330 3350 50080 3365
rect 53285 3405 55035 3420
rect 53285 3365 53300 3405
rect 53340 3365 54980 3405
rect 55020 3365 55035 3405
rect 53285 3350 55035 3365
rect 58240 3405 59990 3420
rect 58240 3365 58255 3405
rect 58295 3365 59935 3405
rect 59975 3365 59990 3405
rect 58240 3350 59990 3365
rect 63195 3405 64945 3420
rect 63195 3365 63210 3405
rect 63250 3365 64890 3405
rect 64930 3365 64945 3405
rect 63195 3350 64945 3365
rect 68150 3405 69900 3420
rect 68150 3365 68165 3405
rect 68205 3365 69845 3405
rect 69885 3365 69900 3405
rect 68150 3350 69900 3365
rect 73105 3405 74855 3420
rect 73105 3365 73120 3405
rect 73160 3365 74800 3405
rect 74840 3365 74855 3405
rect 73105 3350 74855 3365
rect 660 3120 730 3135
rect 660 3080 675 3120
rect 715 3080 730 3120
rect 660 2850 730 3080
rect -175 2835 730 2850
rect -175 2800 675 2835
rect 715 2800 730 2835
rect -175 2785 730 2800
rect -175 1775 -100 2785
rect 660 2490 730 2785
rect 660 2450 675 2490
rect 715 2450 730 2490
rect 660 2435 730 2450
rect 1860 2835 1930 3135
rect 1860 2800 1875 2835
rect 1915 2800 1930 2835
rect 1860 2435 1930 2800
rect 2090 2520 2175 3050
rect 2340 2835 2410 3135
rect 2340 2800 2355 2835
rect 2395 2800 2410 2835
rect 2340 2435 2410 2800
rect 3540 2835 3610 3135
rect 3540 2800 3555 2835
rect 3595 2800 3610 2835
rect 3540 2435 3610 2800
rect 4595 2265 4670 3350
rect 5615 3120 5685 3135
rect 5615 3080 5630 3120
rect 5670 3080 5685 3120
rect 5615 2835 5685 3080
rect 5615 2800 5630 2835
rect 5670 2800 5685 2835
rect 5615 2490 5685 2800
rect 5615 2450 5630 2490
rect 5670 2450 5685 2490
rect 5615 2435 5685 2450
rect 6815 3120 6885 3135
rect 6815 3080 6830 3120
rect 6870 3080 6885 3120
rect 6815 2835 6885 3080
rect 7295 3120 7365 3135
rect 7295 3080 7310 3120
rect 7350 3080 7365 3120
rect 6815 2800 6830 2835
rect 6870 2800 6885 2835
rect 6815 2490 6885 2800
rect 7045 2520 7130 3050
rect 7295 2835 7365 3080
rect 7295 2800 7310 2835
rect 7350 2800 7365 2835
rect 6815 2450 6830 2490
rect 6870 2450 6885 2490
rect 6815 2435 6885 2450
rect 7295 2490 7365 2800
rect 7295 2450 7310 2490
rect 7350 2450 7365 2490
rect 7295 2435 7365 2450
rect 8495 3120 8565 3135
rect 8495 3080 8510 3120
rect 8550 3080 8565 3120
rect 8495 2835 8565 3080
rect 8495 2800 8510 2835
rect 8550 2800 8565 2835
rect 8495 2490 8565 2800
rect 8495 2450 8510 2490
rect 8550 2450 8565 2490
rect 8495 2435 8565 2450
rect 9550 2265 9625 3350
rect 10570 3120 10640 3135
rect 10570 3080 10585 3120
rect 10625 3080 10640 3120
rect 10570 2835 10640 3080
rect 10570 2800 10585 2835
rect 10625 2800 10640 2835
rect 10570 2490 10640 2800
rect 10570 2450 10585 2490
rect 10625 2450 10640 2490
rect 10570 2435 10640 2450
rect 11770 3120 11840 3135
rect 11770 3080 11785 3120
rect 11825 3080 11840 3120
rect 11770 2835 11840 3080
rect 12250 3120 12320 3135
rect 12250 3080 12265 3120
rect 12305 3080 12320 3120
rect 11770 2800 11785 2835
rect 11825 2800 11840 2835
rect 11770 2490 11840 2800
rect 12000 2520 12085 3050
rect 12250 2835 12320 3080
rect 12250 2800 12265 2835
rect 12305 2800 12320 2835
rect 11770 2450 11785 2490
rect 11825 2450 11840 2490
rect 11770 2435 11840 2450
rect 12250 2490 12320 2800
rect 12250 2450 12265 2490
rect 12305 2450 12320 2490
rect 12250 2435 12320 2450
rect 13450 3120 13520 3135
rect 13450 3080 13465 3120
rect 13505 3080 13520 3120
rect 13450 2835 13520 3080
rect 13450 2800 13465 2835
rect 13505 2800 13520 2835
rect 13450 2490 13520 2800
rect 13450 2450 13465 2490
rect 13505 2450 13520 2490
rect 13450 2435 13520 2450
rect 14505 2265 14580 3350
rect 15525 3120 15595 3135
rect 15525 3080 15540 3120
rect 15580 3080 15595 3120
rect 15525 2835 15595 3080
rect 15525 2800 15540 2835
rect 15580 2800 15595 2835
rect 15525 2490 15595 2800
rect 15525 2450 15540 2490
rect 15580 2450 15595 2490
rect 15525 2435 15595 2450
rect 16725 3120 16795 3135
rect 16725 3080 16740 3120
rect 16780 3080 16795 3120
rect 16725 2835 16795 3080
rect 17205 3120 17275 3135
rect 17205 3080 17220 3120
rect 17260 3080 17275 3120
rect 16725 2800 16740 2835
rect 16780 2800 16795 2835
rect 16725 2490 16795 2800
rect 16955 2520 17040 3050
rect 17205 2835 17275 3080
rect 17205 2800 17220 2835
rect 17260 2800 17275 2835
rect 16725 2450 16740 2490
rect 16780 2450 16795 2490
rect 16725 2435 16795 2450
rect 17205 2490 17275 2800
rect 17205 2450 17220 2490
rect 17260 2450 17275 2490
rect 17205 2435 17275 2450
rect 18405 3120 18475 3135
rect 18405 3080 18420 3120
rect 18460 3080 18475 3120
rect 18405 2835 18475 3080
rect 18405 2800 18420 2835
rect 18460 2800 18475 2835
rect 18405 2490 18475 2800
rect 18405 2450 18420 2490
rect 18460 2450 18475 2490
rect 18405 2435 18475 2450
rect 19460 2265 19535 3350
rect 20480 3120 20550 3135
rect 20480 3080 20495 3120
rect 20535 3080 20550 3120
rect 20480 2835 20550 3080
rect 20480 2800 20495 2835
rect 20535 2800 20550 2835
rect 20480 2490 20550 2800
rect 20480 2450 20495 2490
rect 20535 2450 20550 2490
rect 20480 2435 20550 2450
rect 21680 3120 21750 3135
rect 21680 3080 21695 3120
rect 21735 3080 21750 3120
rect 21680 2835 21750 3080
rect 22160 3120 22230 3135
rect 22160 3080 22175 3120
rect 22215 3080 22230 3120
rect 21680 2800 21695 2835
rect 21735 2800 21750 2835
rect 21680 2490 21750 2800
rect 21910 2520 21995 3050
rect 22160 2835 22230 3080
rect 22160 2800 22175 2835
rect 22215 2800 22230 2835
rect 21680 2450 21695 2490
rect 21735 2450 21750 2490
rect 21680 2435 21750 2450
rect 22160 2490 22230 2800
rect 22160 2450 22175 2490
rect 22215 2450 22230 2490
rect 22160 2435 22230 2450
rect 23360 3120 23430 3135
rect 23360 3080 23375 3120
rect 23415 3080 23430 3120
rect 23360 2835 23430 3080
rect 23360 2800 23375 2835
rect 23415 2800 23430 2835
rect 23360 2490 23430 2800
rect 23360 2450 23375 2490
rect 23415 2450 23430 2490
rect 23360 2435 23430 2450
rect 24415 2265 24490 3350
rect 25435 3120 25505 3135
rect 25435 3080 25450 3120
rect 25490 3080 25505 3120
rect 25435 2835 25505 3080
rect 25435 2800 25450 2835
rect 25490 2800 25505 2835
rect 25435 2490 25505 2800
rect 25435 2450 25450 2490
rect 25490 2450 25505 2490
rect 25435 2435 25505 2450
rect 26635 3120 26705 3135
rect 26635 3080 26650 3120
rect 26690 3080 26705 3120
rect 26635 2835 26705 3080
rect 27115 3120 27185 3135
rect 27115 3080 27130 3120
rect 27170 3080 27185 3120
rect 26635 2800 26650 2835
rect 26690 2800 26705 2835
rect 26635 2490 26705 2800
rect 26865 2520 26950 3050
rect 27115 2835 27185 3080
rect 27115 2800 27130 2835
rect 27170 2800 27185 2835
rect 26635 2450 26650 2490
rect 26690 2450 26705 2490
rect 26635 2435 26705 2450
rect 27115 2490 27185 2800
rect 27115 2450 27130 2490
rect 27170 2450 27185 2490
rect 27115 2435 27185 2450
rect 28315 3120 28385 3135
rect 28315 3080 28330 3120
rect 28370 3080 28385 3120
rect 28315 2835 28385 3080
rect 28315 2800 28330 2835
rect 28370 2800 28385 2835
rect 28315 2490 28385 2800
rect 28315 2450 28330 2490
rect 28370 2450 28385 2490
rect 28315 2435 28385 2450
rect 29370 2265 29445 3350
rect 30390 3120 30460 3135
rect 30390 3080 30405 3120
rect 30445 3080 30460 3120
rect 30390 2835 30460 3080
rect 30390 2800 30405 2835
rect 30445 2800 30460 2835
rect 30390 2490 30460 2800
rect 30390 2450 30405 2490
rect 30445 2450 30460 2490
rect 30390 2435 30460 2450
rect 31590 3120 31660 3135
rect 31590 3080 31605 3120
rect 31645 3080 31660 3120
rect 31590 2835 31660 3080
rect 32070 3120 32140 3135
rect 32070 3080 32085 3120
rect 32125 3080 32140 3120
rect 31590 2800 31605 2835
rect 31645 2800 31660 2835
rect 31590 2490 31660 2800
rect 31820 2520 31905 3050
rect 32070 2835 32140 3080
rect 32070 2800 32085 2835
rect 32125 2800 32140 2835
rect 31590 2450 31605 2490
rect 31645 2450 31660 2490
rect 31590 2435 31660 2450
rect 32070 2490 32140 2800
rect 32070 2450 32085 2490
rect 32125 2450 32140 2490
rect 32070 2435 32140 2450
rect 33270 3120 33340 3135
rect 33270 3080 33285 3120
rect 33325 3080 33340 3120
rect 33270 2835 33340 3080
rect 33270 2800 33285 2835
rect 33325 2800 33340 2835
rect 33270 2490 33340 2800
rect 33270 2450 33285 2490
rect 33325 2450 33340 2490
rect 33270 2435 33340 2450
rect 34325 2265 34400 3350
rect 35345 3120 35415 3135
rect 35345 3080 35360 3120
rect 35400 3080 35415 3120
rect 35345 2835 35415 3080
rect 35345 2800 35360 2835
rect 35400 2800 35415 2835
rect 35345 2490 35415 2800
rect 35345 2450 35360 2490
rect 35400 2450 35415 2490
rect 35345 2435 35415 2450
rect 36545 3120 36615 3135
rect 36545 3080 36560 3120
rect 36600 3080 36615 3120
rect 36545 2835 36615 3080
rect 37025 3120 37095 3135
rect 37025 3080 37040 3120
rect 37080 3080 37095 3120
rect 36545 2800 36560 2835
rect 36600 2800 36615 2835
rect 36545 2490 36615 2800
rect 36775 2520 36860 3050
rect 37025 2835 37095 3080
rect 37025 2800 37040 2835
rect 37080 2800 37095 2835
rect 36545 2450 36560 2490
rect 36600 2450 36615 2490
rect 36545 2435 36615 2450
rect 37025 2490 37095 2800
rect 37025 2450 37040 2490
rect 37080 2450 37095 2490
rect 37025 2435 37095 2450
rect 38225 3120 38295 3135
rect 38225 3080 38240 3120
rect 38280 3080 38295 3120
rect 38225 2835 38295 3080
rect 38225 2800 38240 2835
rect 38280 2800 38295 2835
rect 38225 2490 38295 2800
rect 38225 2450 38240 2490
rect 38280 2450 38295 2490
rect 38225 2435 38295 2450
rect 39280 2265 39355 3350
rect 40300 3120 40370 3135
rect 40300 3080 40315 3120
rect 40355 3080 40370 3120
rect 40300 2835 40370 3080
rect 40300 2800 40315 2835
rect 40355 2800 40370 2835
rect 40300 2490 40370 2800
rect 40300 2450 40315 2490
rect 40355 2450 40370 2490
rect 40300 2435 40370 2450
rect 41500 3120 41570 3135
rect 41500 3080 41515 3120
rect 41555 3080 41570 3120
rect 41500 2835 41570 3080
rect 41980 3120 42050 3135
rect 41980 3080 41995 3120
rect 42035 3080 42050 3120
rect 41500 2800 41515 2835
rect 41555 2800 41570 2835
rect 41500 2490 41570 2800
rect 41730 2520 41815 3050
rect 41980 2835 42050 3080
rect 41980 2800 41995 2835
rect 42035 2800 42050 2835
rect 41500 2450 41515 2490
rect 41555 2450 41570 2490
rect 41500 2435 41570 2450
rect 41980 2490 42050 2800
rect 41980 2450 41995 2490
rect 42035 2450 42050 2490
rect 41980 2435 42050 2450
rect 43180 3120 43250 3135
rect 43180 3080 43195 3120
rect 43235 3080 43250 3120
rect 43180 2835 43250 3080
rect 43180 2800 43195 2835
rect 43235 2800 43250 2835
rect 43180 2490 43250 2800
rect 43180 2450 43195 2490
rect 43235 2450 43250 2490
rect 43180 2435 43250 2450
rect 44235 2265 44310 3350
rect 45255 3120 45325 3135
rect 45255 3080 45270 3120
rect 45310 3080 45325 3120
rect 45255 2835 45325 3080
rect 45255 2800 45270 2835
rect 45310 2800 45325 2835
rect 45255 2490 45325 2800
rect 45255 2450 45270 2490
rect 45310 2450 45325 2490
rect 45255 2435 45325 2450
rect 46455 3120 46525 3135
rect 46455 3080 46470 3120
rect 46510 3080 46525 3120
rect 46455 2835 46525 3080
rect 46935 3120 47005 3135
rect 46935 3080 46950 3120
rect 46990 3080 47005 3120
rect 46455 2800 46470 2835
rect 46510 2800 46525 2835
rect 46455 2490 46525 2800
rect 46685 2520 46770 3050
rect 46935 2835 47005 3080
rect 46935 2800 46950 2835
rect 46990 2800 47005 2835
rect 46455 2450 46470 2490
rect 46510 2450 46525 2490
rect 46455 2435 46525 2450
rect 46935 2490 47005 2800
rect 46935 2450 46950 2490
rect 46990 2450 47005 2490
rect 46935 2435 47005 2450
rect 48135 3120 48205 3135
rect 48135 3080 48150 3120
rect 48190 3080 48205 3120
rect 48135 2835 48205 3080
rect 48135 2800 48150 2835
rect 48190 2800 48205 2835
rect 48135 2490 48205 2800
rect 48135 2450 48150 2490
rect 48190 2450 48205 2490
rect 48135 2435 48205 2450
rect 49190 2265 49265 3350
rect 50210 3120 50280 3135
rect 50210 3080 50225 3120
rect 50265 3080 50280 3120
rect 50210 2835 50280 3080
rect 50210 2800 50225 2835
rect 50265 2800 50280 2835
rect 50210 2490 50280 2800
rect 50210 2450 50225 2490
rect 50265 2450 50280 2490
rect 50210 2435 50280 2450
rect 51410 3120 51480 3135
rect 51410 3080 51425 3120
rect 51465 3080 51480 3120
rect 51410 2835 51480 3080
rect 51890 3120 51960 3135
rect 51890 3080 51905 3120
rect 51945 3080 51960 3120
rect 51410 2800 51425 2835
rect 51465 2800 51480 2835
rect 51410 2490 51480 2800
rect 51640 2520 51725 3050
rect 51890 2835 51960 3080
rect 51890 2800 51905 2835
rect 51945 2800 51960 2835
rect 51410 2450 51425 2490
rect 51465 2450 51480 2490
rect 51410 2435 51480 2450
rect 51890 2490 51960 2800
rect 51890 2450 51905 2490
rect 51945 2450 51960 2490
rect 51890 2435 51960 2450
rect 53090 3120 53160 3135
rect 53090 3080 53105 3120
rect 53145 3080 53160 3120
rect 53090 2835 53160 3080
rect 53090 2800 53105 2835
rect 53145 2800 53160 2835
rect 53090 2490 53160 2800
rect 53090 2450 53105 2490
rect 53145 2450 53160 2490
rect 53090 2435 53160 2450
rect 54145 2265 54220 3350
rect 55165 3120 55235 3135
rect 55165 3080 55180 3120
rect 55220 3080 55235 3120
rect 55165 2835 55235 3080
rect 55165 2800 55180 2835
rect 55220 2800 55235 2835
rect 55165 2490 55235 2800
rect 55165 2450 55180 2490
rect 55220 2450 55235 2490
rect 55165 2435 55235 2450
rect 56365 3120 56435 3135
rect 56365 3080 56380 3120
rect 56420 3080 56435 3120
rect 56365 2835 56435 3080
rect 56845 3120 56915 3135
rect 56845 3080 56860 3120
rect 56900 3080 56915 3120
rect 56365 2800 56380 2835
rect 56420 2800 56435 2835
rect 56365 2490 56435 2800
rect 56595 2520 56680 3050
rect 56845 2835 56915 3080
rect 56845 2800 56860 2835
rect 56900 2800 56915 2835
rect 56365 2450 56380 2490
rect 56420 2450 56435 2490
rect 56365 2435 56435 2450
rect 56845 2490 56915 2800
rect 56845 2450 56860 2490
rect 56900 2450 56915 2490
rect 56845 2435 56915 2450
rect 58045 3120 58115 3135
rect 58045 3080 58060 3120
rect 58100 3080 58115 3120
rect 58045 2835 58115 3080
rect 58045 2800 58060 2835
rect 58100 2800 58115 2835
rect 58045 2490 58115 2800
rect 58045 2450 58060 2490
rect 58100 2450 58115 2490
rect 58045 2435 58115 2450
rect 59100 2265 59175 3350
rect 60120 3120 60190 3135
rect 60120 3080 60135 3120
rect 60175 3080 60190 3120
rect 60120 2835 60190 3080
rect 60120 2800 60135 2835
rect 60175 2800 60190 2835
rect 60120 2490 60190 2800
rect 60120 2450 60135 2490
rect 60175 2450 60190 2490
rect 60120 2435 60190 2450
rect 61320 3120 61390 3135
rect 61320 3080 61335 3120
rect 61375 3080 61390 3120
rect 61320 2835 61390 3080
rect 61800 3120 61870 3135
rect 61800 3080 61815 3120
rect 61855 3080 61870 3120
rect 61320 2800 61335 2835
rect 61375 2800 61390 2835
rect 61320 2490 61390 2800
rect 61550 2520 61635 3050
rect 61800 2835 61870 3080
rect 61800 2800 61815 2835
rect 61855 2800 61870 2835
rect 61320 2450 61335 2490
rect 61375 2450 61390 2490
rect 61320 2435 61390 2450
rect 61800 2490 61870 2800
rect 61800 2450 61815 2490
rect 61855 2450 61870 2490
rect 61800 2435 61870 2450
rect 63000 3120 63070 3135
rect 63000 3080 63015 3120
rect 63055 3080 63070 3120
rect 63000 2835 63070 3080
rect 63000 2800 63015 2835
rect 63055 2800 63070 2835
rect 63000 2490 63070 2800
rect 63000 2450 63015 2490
rect 63055 2450 63070 2490
rect 63000 2435 63070 2450
rect 64055 2265 64130 3350
rect 65075 3120 65145 3135
rect 65075 3080 65090 3120
rect 65130 3080 65145 3120
rect 65075 2835 65145 3080
rect 65075 2800 65090 2835
rect 65130 2800 65145 2835
rect 65075 2490 65145 2800
rect 65075 2450 65090 2490
rect 65130 2450 65145 2490
rect 65075 2435 65145 2450
rect 66275 3120 66345 3135
rect 66275 3080 66290 3120
rect 66330 3080 66345 3120
rect 66275 2835 66345 3080
rect 66755 3120 66825 3135
rect 66755 3080 66770 3120
rect 66810 3080 66825 3120
rect 66275 2800 66290 2835
rect 66330 2800 66345 2835
rect 66275 2490 66345 2800
rect 66505 2520 66590 3050
rect 66755 2835 66825 3080
rect 66755 2800 66770 2835
rect 66810 2800 66825 2835
rect 66275 2450 66290 2490
rect 66330 2450 66345 2490
rect 66275 2435 66345 2450
rect 66755 2490 66825 2800
rect 66755 2450 66770 2490
rect 66810 2450 66825 2490
rect 66755 2435 66825 2450
rect 67955 3120 68025 3135
rect 67955 3080 67970 3120
rect 68010 3080 68025 3120
rect 67955 2835 68025 3080
rect 67955 2800 67970 2835
rect 68010 2800 68025 2835
rect 67955 2490 68025 2800
rect 67955 2450 67970 2490
rect 68010 2450 68025 2490
rect 67955 2435 68025 2450
rect 69010 2265 69085 3350
rect 70030 3120 70100 3135
rect 70030 3080 70045 3120
rect 70085 3080 70100 3120
rect 70030 2835 70100 3080
rect 70030 2800 70045 2835
rect 70085 2800 70100 2835
rect 70030 2490 70100 2800
rect 70030 2450 70045 2490
rect 70085 2450 70100 2490
rect 70030 2435 70100 2450
rect 71230 3120 71300 3135
rect 71230 3080 71245 3120
rect 71285 3080 71300 3120
rect 71230 2835 71300 3080
rect 71710 3120 71780 3135
rect 71710 3080 71725 3120
rect 71765 3080 71780 3120
rect 71230 2800 71245 2835
rect 71285 2800 71300 2835
rect 71230 2490 71300 2800
rect 71460 2520 71545 3050
rect 71710 2835 71780 3080
rect 71710 2800 71725 2835
rect 71765 2800 71780 2835
rect 71230 2450 71245 2490
rect 71285 2450 71300 2490
rect 71230 2435 71300 2450
rect 71710 2490 71780 2800
rect 71710 2450 71725 2490
rect 71765 2450 71780 2490
rect 71710 2435 71780 2450
rect 72910 3120 72980 3135
rect 72910 3080 72925 3120
rect 72965 3080 72980 3120
rect 72910 2835 72980 3080
rect 72910 2800 72925 2835
rect 72965 2800 72980 2835
rect 72910 2490 72980 2800
rect 72910 2450 72925 2490
rect 72965 2450 72980 2490
rect 72910 2435 72980 2450
rect 73965 2265 74040 3350
rect 74985 3120 75055 3135
rect 74985 3080 75000 3120
rect 75040 3080 75055 3120
rect 74985 2835 75055 3080
rect 74985 2800 75000 2835
rect 75040 2800 75055 2835
rect 74985 2490 75055 2800
rect 74985 2450 75000 2490
rect 75040 2450 75055 2490
rect 74985 2435 75055 2450
rect 76185 3120 76255 3135
rect 76185 3080 76200 3120
rect 76240 3080 76255 3120
rect 76185 2835 76255 3080
rect 76665 3120 76735 3135
rect 76665 3080 76680 3120
rect 76720 3080 76735 3120
rect 76185 2800 76200 2835
rect 76240 2800 76255 2835
rect 76185 2490 76255 2800
rect 76415 2520 76500 3050
rect 76665 2835 76735 3080
rect 76665 2800 76680 2835
rect 76720 2800 76735 2835
rect 76185 2450 76200 2490
rect 76240 2450 76255 2490
rect 76185 2435 76255 2450
rect 76665 2490 76735 2800
rect 76665 2450 76680 2490
rect 76720 2450 76735 2490
rect 76665 2435 76735 2450
rect 77865 3120 77935 3135
rect 77865 3080 77880 3120
rect 77920 3080 77935 3120
rect 77865 2835 77935 3080
rect 77865 2800 77880 2835
rect 77920 2800 77935 2835
rect 77865 2490 77935 2800
rect 77865 2450 77880 2490
rect 77920 2450 77935 2490
rect 77865 2435 77935 2450
rect 3735 2195 5485 2265
rect 8690 2250 10440 2265
rect 8690 2210 8705 2250
rect 8745 2210 10385 2250
rect 10425 2210 10440 2250
rect 8690 2195 10440 2210
rect 13645 2250 15395 2265
rect 13645 2210 13660 2250
rect 13700 2210 15340 2250
rect 15380 2210 15395 2250
rect 13645 2195 15395 2210
rect 18600 2250 20350 2265
rect 18600 2210 18615 2250
rect 18655 2210 20295 2250
rect 20335 2210 20350 2250
rect 18600 2195 20350 2210
rect 23555 2250 25305 2265
rect 23555 2210 23570 2250
rect 23610 2210 25250 2250
rect 25290 2210 25305 2250
rect 23555 2195 25305 2210
rect 28510 2250 30260 2265
rect 28510 2210 28525 2250
rect 28565 2210 30205 2250
rect 30245 2210 30260 2250
rect 28510 2195 30260 2210
rect 33465 2250 35215 2265
rect 33465 2210 33480 2250
rect 33520 2210 35160 2250
rect 35200 2210 35215 2250
rect 33465 2195 35215 2210
rect 38420 2250 40170 2265
rect 38420 2210 38435 2250
rect 38475 2210 40115 2250
rect 40155 2210 40170 2250
rect 38420 2195 40170 2210
rect 43375 2250 45125 2265
rect 43375 2210 43390 2250
rect 43430 2210 45070 2250
rect 45110 2210 45125 2250
rect 43375 2195 45125 2210
rect 48330 2250 50080 2265
rect 48330 2210 48345 2250
rect 48385 2210 50025 2250
rect 50065 2210 50080 2250
rect 48330 2195 50080 2210
rect 53285 2250 55035 2265
rect 53285 2210 53300 2250
rect 53340 2210 54980 2250
rect 55020 2210 55035 2250
rect 53285 2195 55035 2210
rect 58240 2250 59990 2265
rect 58240 2210 58255 2250
rect 58295 2210 59935 2250
rect 59975 2210 59990 2250
rect 58240 2195 59990 2210
rect 63195 2250 64945 2265
rect 63195 2210 63210 2250
rect 63250 2210 64890 2250
rect 64930 2210 64945 2250
rect 63195 2195 64945 2210
rect 68150 2250 69900 2265
rect 68150 2210 68165 2250
rect 68205 2210 69845 2250
rect 69885 2210 69900 2250
rect 68150 2195 69900 2210
rect 73105 2250 74855 2265
rect 73105 2210 73120 2250
rect 73160 2210 74800 2250
rect 74840 2210 74855 2250
rect 73105 2195 74855 2210
rect -345 1700 -100 1775
rect 4595 345 4670 2195
rect 9550 345 9625 2195
rect 14505 345 14580 2195
rect 19460 345 19535 2195
rect 24415 345 24490 2195
rect 29370 345 29445 2195
rect 34325 345 34400 2195
rect 39280 345 39355 2195
rect 44235 345 44310 2195
rect 49190 345 49265 2195
rect 54145 345 54220 2195
rect 59100 345 59175 2195
rect 64055 345 64130 2195
rect 69010 345 69085 2195
rect 73965 345 74040 2195
rect 3735 275 5485 345
rect 8690 330 10440 345
rect 8690 290 8705 330
rect 8745 290 10385 330
rect 10425 290 10440 330
rect 8690 275 10440 290
rect 13645 330 15395 345
rect 13645 290 13660 330
rect 13700 290 15340 330
rect 15380 290 15395 330
rect 13645 275 15395 290
rect 18600 330 20350 345
rect 18600 290 18615 330
rect 18655 290 20295 330
rect 20335 290 20350 330
rect 18600 275 20350 290
rect 23555 330 25305 345
rect 23555 290 23570 330
rect 23610 290 25250 330
rect 25290 290 25305 330
rect 23555 275 25305 290
rect 28510 330 30260 345
rect 28510 290 28525 330
rect 28565 290 30205 330
rect 30245 290 30260 330
rect 28510 275 30260 290
rect 33465 330 35215 345
rect 33465 290 33480 330
rect 33520 290 35160 330
rect 35200 290 35215 330
rect 33465 275 35215 290
rect 38420 330 40170 345
rect 38420 290 38435 330
rect 38475 290 40115 330
rect 40155 290 40170 330
rect 38420 275 40170 290
rect 43375 330 45125 345
rect 43375 290 43390 330
rect 43430 290 45070 330
rect 45110 290 45125 330
rect 43375 275 45125 290
rect 48330 330 50080 345
rect 48330 290 48345 330
rect 48385 290 50025 330
rect 50065 290 50080 330
rect 48330 275 50080 290
rect 53285 330 55035 345
rect 53285 290 53300 330
rect 53340 290 54980 330
rect 55020 290 55035 330
rect 53285 275 55035 290
rect 58240 330 59990 345
rect 58240 290 58255 330
rect 58295 290 59935 330
rect 59975 290 59990 330
rect 58240 275 59990 290
rect 63195 330 64945 345
rect 63195 290 63210 330
rect 63250 290 64890 330
rect 64930 290 64945 330
rect 63195 275 64945 290
rect 68150 330 69900 345
rect 68150 290 68165 330
rect 68205 290 69845 330
rect 69885 290 69900 330
rect 68150 275 69900 290
rect 73105 330 74855 345
rect 73105 290 73120 330
rect 73160 290 74800 330
rect 74840 290 74855 330
rect 73105 275 74855 290
rect 2090 -265 2175 55
rect 7045 40 7130 55
rect 7045 -10 7060 40
rect 7115 -10 7130 40
rect 7045 -265 7130 -10
rect 12000 40 12085 55
rect 12000 -10 12015 40
rect 12070 -10 12085 40
rect 12000 -265 12085 -10
rect 16955 40 17040 55
rect 16955 -10 16970 40
rect 17025 -10 17040 40
rect 16955 -265 17040 -10
rect 21910 40 21995 55
rect 21910 -10 21925 40
rect 21980 -10 21995 40
rect 21910 -265 21995 -10
rect 26865 40 26950 55
rect 26865 -10 26880 40
rect 26935 -10 26950 40
rect 26865 -265 26950 -10
rect 31820 40 31905 55
rect 31820 -10 31835 40
rect 31890 -10 31905 40
rect 31820 -265 31905 -10
rect 36775 40 36860 55
rect 36775 -10 36790 40
rect 36845 -10 36860 40
rect 36775 -265 36860 -10
rect 41730 40 41815 55
rect 41730 -10 41745 40
rect 41800 -10 41815 40
rect 41730 -265 41815 -10
rect 46685 40 46770 55
rect 46685 -10 46700 40
rect 46755 -10 46770 40
rect 46685 -265 46770 -10
rect 51640 40 51725 55
rect 51640 -10 51655 40
rect 51710 -10 51725 40
rect 51640 -265 51725 -10
rect 56595 40 56680 55
rect 56595 -10 56610 40
rect 56665 -10 56680 40
rect 56595 -265 56680 -10
rect 61550 40 61635 55
rect 61550 -10 61565 40
rect 61620 -10 61635 40
rect 61550 -265 61635 -10
rect 66505 40 66590 55
rect 66505 -10 66520 40
rect 66575 -10 66590 40
rect 66505 -265 66590 -10
rect 71460 40 71545 55
rect 71460 -10 71475 40
rect 71530 -10 71545 40
rect 71460 -265 71545 -10
rect 76415 40 76500 55
rect 76415 -10 76430 40
rect 76485 -10 76500 40
rect 76415 -265 76500 -10
rect 78745 -265 78830 11985
rect 2090 -345 78830 -265
<< viali >>
rect -330 11920 -200 12050
rect 8705 11435 8745 11475
rect 10385 11435 10425 11475
rect 13660 11435 13700 11475
rect 15340 11435 15380 11475
rect 18615 11435 18655 11475
rect 20295 11435 20335 11475
rect 23570 11435 23610 11475
rect 25250 11435 25290 11475
rect 28525 11435 28565 11475
rect 30205 11435 30245 11475
rect 33480 11435 33520 11475
rect 35160 11435 35200 11475
rect 38435 11435 38475 11475
rect 40115 11435 40155 11475
rect 43390 11435 43430 11475
rect 45070 11435 45110 11475
rect 48345 11435 48385 11475
rect 50025 11435 50065 11475
rect 53300 11435 53340 11475
rect 54980 11435 55020 11475
rect 58255 11435 58295 11475
rect 59935 11435 59975 11475
rect 63210 11435 63250 11475
rect 64890 11435 64930 11475
rect 68165 11435 68205 11475
rect 69845 11435 69885 11475
rect 73120 11435 73160 11475
rect 74800 11435 74840 11475
rect 8705 9515 8745 9555
rect 10385 9515 10425 9555
rect 13660 9515 13700 9555
rect 15340 9515 15380 9555
rect 18615 9515 18655 9555
rect 20295 9515 20335 9555
rect 23570 9515 23610 9555
rect 25250 9515 25290 9555
rect 28525 9515 28565 9555
rect 30205 9515 30245 9555
rect 33480 9515 33520 9555
rect 35160 9515 35200 9555
rect 38435 9515 38475 9555
rect 40115 9515 40155 9555
rect 43390 9515 43430 9555
rect 45070 9515 45110 9555
rect 48345 9515 48385 9555
rect 50025 9515 50065 9555
rect 53300 9515 53340 9555
rect 54980 9515 55020 9555
rect 58255 9515 58295 9555
rect 59935 9515 59975 9555
rect 63210 9515 63250 9555
rect 64890 9515 64930 9555
rect 68165 9515 68205 9555
rect 69845 9515 69885 9555
rect 73120 9515 73160 9555
rect 74800 9515 74840 9555
rect 675 8900 715 8935
rect 1875 8900 1915 8935
rect 2355 8900 2395 8935
rect 3555 8900 3595 8935
rect 5630 9230 5670 9270
rect 5630 8900 5670 8935
rect 5630 8600 5670 8640
rect 6830 9230 6870 9270
rect 7310 9230 7350 9270
rect 6830 8900 6870 8935
rect 7310 8900 7350 8935
rect 6830 8600 6870 8640
rect 7310 8600 7350 8640
rect 8510 9230 8550 9270
rect 8510 8900 8550 8935
rect 8510 8600 8550 8640
rect 10585 9230 10625 9270
rect 10585 8900 10625 8935
rect 10585 8600 10625 8640
rect 11785 9230 11825 9270
rect 12265 9230 12305 9270
rect 11785 8900 11825 8935
rect 12265 8900 12305 8935
rect 11785 8600 11825 8640
rect 12265 8600 12305 8640
rect 13465 9230 13505 9270
rect 13465 8900 13505 8935
rect 13465 8600 13505 8640
rect 15540 9230 15580 9270
rect 15540 8900 15580 8935
rect 15540 8600 15580 8640
rect 16740 9230 16780 9270
rect 17220 9230 17260 9270
rect 16740 8900 16780 8935
rect 17220 8900 17260 8935
rect 16740 8600 16780 8640
rect 17220 8600 17260 8640
rect 18420 9230 18460 9270
rect 18420 8900 18460 8935
rect 18420 8600 18460 8640
rect 20495 9230 20535 9270
rect 20495 8900 20535 8935
rect 20495 8600 20535 8640
rect 21695 9230 21735 9270
rect 22175 9230 22215 9270
rect 21695 8900 21735 8935
rect 22175 8900 22215 8935
rect 21695 8600 21735 8640
rect 22175 8600 22215 8640
rect 23375 9230 23415 9270
rect 23375 8900 23415 8935
rect 23375 8600 23415 8640
rect 25450 9230 25490 9270
rect 25450 8900 25490 8935
rect 25450 8600 25490 8640
rect 26650 9230 26690 9270
rect 27130 9230 27170 9270
rect 26650 8900 26690 8935
rect 27130 8900 27170 8935
rect 26650 8600 26690 8640
rect 27130 8600 27170 8640
rect 28330 9230 28370 9270
rect 28330 8900 28370 8935
rect 28330 8600 28370 8640
rect 30405 9230 30445 9270
rect 30405 8900 30445 8935
rect 30405 8600 30445 8640
rect 31605 9230 31645 9270
rect 32085 9230 32125 9270
rect 31605 8900 31645 8935
rect 32085 8900 32125 8935
rect 31605 8600 31645 8640
rect 32085 8600 32125 8640
rect 33285 9230 33325 9270
rect 33285 8900 33325 8935
rect 33285 8600 33325 8640
rect 35360 9230 35400 9270
rect 35360 8900 35400 8935
rect 35360 8600 35400 8640
rect 36560 9230 36600 9270
rect 37040 9230 37080 9270
rect 36560 8900 36600 8935
rect 37040 8900 37080 8935
rect 36560 8600 36600 8640
rect 37040 8600 37080 8640
rect 38240 9230 38280 9270
rect 38240 8900 38280 8935
rect 38240 8600 38280 8640
rect 40315 9230 40355 9270
rect 40315 8900 40355 8935
rect 40315 8600 40355 8640
rect 41515 9230 41555 9270
rect 41995 9230 42035 9270
rect 41515 8900 41555 8935
rect 41995 8900 42035 8935
rect 41515 8600 41555 8640
rect 41995 8600 42035 8640
rect 43195 9230 43235 9270
rect 43195 8900 43235 8935
rect 43195 8600 43235 8640
rect 45270 9230 45310 9270
rect 45270 8900 45310 8935
rect 45270 8600 45310 8640
rect 46470 9230 46510 9270
rect 46950 9230 46990 9270
rect 46470 8900 46510 8935
rect 46950 8900 46990 8935
rect 46470 8600 46510 8640
rect 46950 8600 46990 8640
rect 48150 9230 48190 9270
rect 48150 8900 48190 8935
rect 48150 8600 48190 8640
rect 50225 9230 50265 9270
rect 50225 8900 50265 8935
rect 50225 8600 50265 8640
rect 51425 9230 51465 9270
rect 51905 9230 51945 9270
rect 51425 8900 51465 8935
rect 51905 8900 51945 8935
rect 51425 8600 51465 8640
rect 51905 8600 51945 8640
rect 53105 9230 53145 9270
rect 53105 8900 53145 8935
rect 53105 8600 53145 8640
rect 55180 9230 55220 9270
rect 55180 8900 55220 8935
rect 55180 8600 55220 8640
rect 56380 9230 56420 9270
rect 56860 9230 56900 9270
rect 56380 8900 56420 8935
rect 56860 8900 56900 8935
rect 56380 8600 56420 8640
rect 56860 8600 56900 8640
rect 58060 9230 58100 9270
rect 58060 8900 58100 8935
rect 58060 8600 58100 8640
rect 60135 9230 60175 9270
rect 60135 8900 60175 8935
rect 60135 8600 60175 8640
rect 61335 9230 61375 9270
rect 61815 9230 61855 9270
rect 61335 8900 61375 8935
rect 61815 8900 61855 8935
rect 61335 8600 61375 8640
rect 61815 8600 61855 8640
rect 63015 9230 63055 9270
rect 63015 8900 63055 8935
rect 63015 8600 63055 8640
rect 65090 9230 65130 9270
rect 65090 8900 65130 8935
rect 65090 8600 65130 8640
rect 66290 9230 66330 9270
rect 66770 9230 66810 9270
rect 66290 8900 66330 8935
rect 66770 8900 66810 8935
rect 66290 8600 66330 8640
rect 66770 8600 66810 8640
rect 67970 9230 68010 9270
rect 67970 8900 68010 8935
rect 67970 8600 68010 8640
rect 70045 9230 70085 9270
rect 70045 8900 70085 8935
rect 70045 8600 70085 8640
rect 71245 9230 71285 9270
rect 71725 9230 71765 9270
rect 71245 8900 71285 8935
rect 71725 8900 71765 8935
rect 71245 8600 71285 8640
rect 71725 8600 71765 8640
rect 72925 9230 72965 9270
rect 72925 8900 72965 8935
rect 72925 8600 72965 8640
rect 75000 9230 75040 9270
rect 75000 8900 75040 8935
rect 75000 8600 75040 8640
rect 76200 9230 76240 9270
rect 76680 9230 76720 9270
rect 76200 8900 76240 8935
rect 76680 8900 76720 8935
rect 76200 8600 76240 8640
rect 76680 8600 76720 8640
rect 77880 9230 77920 9270
rect 77880 8900 77920 8935
rect 77880 8600 77920 8640
rect 8705 8360 8745 8400
rect 10385 8360 10425 8400
rect 13660 8360 13700 8400
rect 15340 8360 15380 8400
rect 18615 8360 18655 8400
rect 20295 8360 20335 8400
rect 23570 8360 23610 8400
rect 25250 8360 25290 8400
rect 28525 8360 28565 8400
rect 30205 8360 30245 8400
rect 33480 8360 33520 8400
rect 35160 8360 35200 8400
rect 38435 8360 38475 8400
rect 40115 8360 40155 8400
rect 43390 8360 43430 8400
rect 45070 8360 45110 8400
rect 48345 8360 48385 8400
rect 50025 8360 50065 8400
rect 53300 8360 53340 8400
rect 54980 8360 55020 8400
rect 58255 8360 58295 8400
rect 59935 8360 59975 8400
rect 63210 8360 63250 8400
rect 64890 8360 64930 8400
rect 68165 8360 68205 8400
rect 69845 8360 69885 8400
rect 73120 8360 73160 8400
rect 74800 8360 74840 8400
rect 8705 6440 8745 6480
rect 10385 6440 10425 6480
rect 13660 6440 13700 6480
rect 15340 6440 15380 6480
rect 18615 6440 18655 6480
rect 20295 6440 20335 6480
rect 23570 6440 23610 6480
rect 25250 6440 25290 6480
rect 28525 6440 28565 6480
rect 30205 6440 30245 6480
rect 33480 6440 33520 6480
rect 35160 6440 35200 6480
rect 38435 6440 38475 6480
rect 40115 6440 40155 6480
rect 43390 6440 43430 6480
rect 45070 6440 45110 6480
rect 48345 6440 48385 6480
rect 50025 6440 50065 6480
rect 53300 6440 53340 6480
rect 54980 6440 55020 6480
rect 58255 6440 58295 6480
rect 59935 6440 59975 6480
rect 63210 6440 63250 6480
rect 64890 6440 64930 6480
rect 68165 6440 68205 6480
rect 69845 6440 69885 6480
rect 73120 6440 73160 6480
rect 74800 6440 74840 6480
rect 675 5850 715 5885
rect 1875 5850 1915 5885
rect 2355 5850 2395 5885
rect 3555 5850 3595 5885
rect 5630 6155 5670 6195
rect 5630 5850 5670 5885
rect 5630 5525 5670 5565
rect 6830 6155 6870 6195
rect 7310 6155 7350 6195
rect 6830 5850 6870 5885
rect 7310 5850 7350 5885
rect 6830 5525 6870 5565
rect 7310 5525 7350 5565
rect 8510 6155 8550 6195
rect 8510 5850 8550 5885
rect 8510 5525 8550 5565
rect 10585 6155 10625 6195
rect 10585 5850 10625 5885
rect 10585 5525 10625 5565
rect 11785 6155 11825 6195
rect 12265 6155 12305 6195
rect 11785 5850 11825 5885
rect 12265 5850 12305 5885
rect 11785 5525 11825 5565
rect 12265 5525 12305 5565
rect 13465 6155 13505 6195
rect 13465 5850 13505 5885
rect 13465 5525 13505 5565
rect 15540 6155 15580 6195
rect 15540 5850 15580 5885
rect 15540 5525 15580 5565
rect 16740 6155 16780 6195
rect 17220 6155 17260 6195
rect 16740 5850 16780 5885
rect 17220 5850 17260 5885
rect 16740 5525 16780 5565
rect 17220 5525 17260 5565
rect 18420 6155 18460 6195
rect 18420 5850 18460 5885
rect 18420 5525 18460 5565
rect 20495 6155 20535 6195
rect 20495 5850 20535 5885
rect 20495 5525 20535 5565
rect 21695 6155 21735 6195
rect 22175 6155 22215 6195
rect 21695 5850 21735 5885
rect 22175 5850 22215 5885
rect 21695 5525 21735 5565
rect 22175 5525 22215 5565
rect 23375 6155 23415 6195
rect 23375 5850 23415 5885
rect 23375 5525 23415 5565
rect 25450 6155 25490 6195
rect 25450 5850 25490 5885
rect 25450 5525 25490 5565
rect 26650 6155 26690 6195
rect 27130 6155 27170 6195
rect 26650 5850 26690 5885
rect 27130 5850 27170 5885
rect 26650 5525 26690 5565
rect 27130 5525 27170 5565
rect 28330 6155 28370 6195
rect 28330 5850 28370 5885
rect 28330 5525 28370 5565
rect 30405 6155 30445 6195
rect 30405 5850 30445 5885
rect 30405 5525 30445 5565
rect 31605 6155 31645 6195
rect 32085 6155 32125 6195
rect 31605 5850 31645 5885
rect 32085 5850 32125 5885
rect 31605 5525 31645 5565
rect 32085 5525 32125 5565
rect 33285 6155 33325 6195
rect 33285 5850 33325 5885
rect 33285 5525 33325 5565
rect 35360 6155 35400 6195
rect 35360 5850 35400 5885
rect 35360 5525 35400 5565
rect 36560 6155 36600 6195
rect 37040 6155 37080 6195
rect 36560 5850 36600 5885
rect 37040 5850 37080 5885
rect 36560 5525 36600 5565
rect 37040 5525 37080 5565
rect 38240 6155 38280 6195
rect 38240 5850 38280 5885
rect 38240 5525 38280 5565
rect 40315 6155 40355 6195
rect 40315 5850 40355 5885
rect 40315 5525 40355 5565
rect 41515 6155 41555 6195
rect 41995 6155 42035 6195
rect 41515 5850 41555 5885
rect 41995 5850 42035 5885
rect 41515 5525 41555 5565
rect 41995 5525 42035 5565
rect 43195 6155 43235 6195
rect 43195 5850 43235 5885
rect 43195 5525 43235 5565
rect 45270 6155 45310 6195
rect 45270 5850 45310 5885
rect 45270 5525 45310 5565
rect 46470 6155 46510 6195
rect 46950 6155 46990 6195
rect 46470 5850 46510 5885
rect 46950 5850 46990 5885
rect 46470 5525 46510 5565
rect 46950 5525 46990 5565
rect 48150 6155 48190 6195
rect 48150 5850 48190 5885
rect 48150 5525 48190 5565
rect 50225 6155 50265 6195
rect 50225 5850 50265 5885
rect 50225 5525 50265 5565
rect 51425 6155 51465 6195
rect 51905 6155 51945 6195
rect 51425 5850 51465 5885
rect 51905 5850 51945 5885
rect 51425 5525 51465 5565
rect 51905 5525 51945 5565
rect 53105 6155 53145 6195
rect 53105 5850 53145 5885
rect 53105 5525 53145 5565
rect 55180 6155 55220 6195
rect 55180 5850 55220 5885
rect 55180 5525 55220 5565
rect 56380 6155 56420 6195
rect 56860 6155 56900 6195
rect 56380 5850 56420 5885
rect 56860 5850 56900 5885
rect 56380 5525 56420 5565
rect 56860 5525 56900 5565
rect 58060 6155 58100 6195
rect 58060 5850 58100 5885
rect 58060 5525 58100 5565
rect 60135 6155 60175 6195
rect 60135 5850 60175 5885
rect 60135 5525 60175 5565
rect 61335 6155 61375 6195
rect 61815 6155 61855 6195
rect 61335 5850 61375 5885
rect 61815 5850 61855 5885
rect 61335 5525 61375 5565
rect 61815 5525 61855 5565
rect 63015 6155 63055 6195
rect 63015 5850 63055 5885
rect 63015 5525 63055 5565
rect 65090 6155 65130 6195
rect 65090 5850 65130 5885
rect 65090 5525 65130 5565
rect 66290 6155 66330 6195
rect 66770 6155 66810 6195
rect 66290 5850 66330 5885
rect 66770 5850 66810 5885
rect 66290 5525 66330 5565
rect 66770 5525 66810 5565
rect 67970 6155 68010 6195
rect 67970 5850 68010 5885
rect 67970 5525 68010 5565
rect 70045 6155 70085 6195
rect 70045 5850 70085 5885
rect 70045 5525 70085 5565
rect 71245 6155 71285 6195
rect 71725 6155 71765 6195
rect 71245 5850 71285 5885
rect 71725 5850 71765 5885
rect 71245 5525 71285 5565
rect 71725 5525 71765 5565
rect 72925 6155 72965 6195
rect 72925 5850 72965 5885
rect 72925 5525 72965 5565
rect 75000 6155 75040 6195
rect 75000 5850 75040 5885
rect 75000 5525 75040 5565
rect 76200 6155 76240 6195
rect 76680 6155 76720 6195
rect 76200 5850 76240 5885
rect 76680 5850 76720 5885
rect 76200 5525 76240 5565
rect 76680 5525 76720 5565
rect 77880 6155 77920 6195
rect 77880 5850 77920 5885
rect 77880 5525 77920 5565
rect 8705 5285 8745 5325
rect 10385 5285 10425 5325
rect 13660 5285 13700 5325
rect 15340 5285 15380 5325
rect 18615 5285 18655 5325
rect 20295 5285 20335 5325
rect 23570 5285 23610 5325
rect 25250 5285 25290 5325
rect 28525 5285 28565 5325
rect 30205 5285 30245 5325
rect 33480 5285 33520 5325
rect 35160 5285 35200 5325
rect 38435 5285 38475 5325
rect 40115 5285 40155 5325
rect 43390 5285 43430 5325
rect 45070 5285 45110 5325
rect 48345 5285 48385 5325
rect 50025 5285 50065 5325
rect 53300 5285 53340 5325
rect 54980 5285 55020 5325
rect 58255 5285 58295 5325
rect 59935 5285 59975 5325
rect 63210 5285 63250 5325
rect 64890 5285 64930 5325
rect 68165 5285 68205 5325
rect 69845 5285 69885 5325
rect 73120 5285 73160 5325
rect 74800 5285 74840 5325
rect 8705 3365 8745 3405
rect 10385 3365 10425 3405
rect 13660 3365 13700 3405
rect 15340 3365 15380 3405
rect 18615 3365 18655 3405
rect 20295 3365 20335 3405
rect 23570 3365 23610 3405
rect 25250 3365 25290 3405
rect 28525 3365 28565 3405
rect 30205 3365 30245 3405
rect 33480 3365 33520 3405
rect 35160 3365 35200 3405
rect 38435 3365 38475 3405
rect 40115 3365 40155 3405
rect 43390 3365 43430 3405
rect 45070 3365 45110 3405
rect 48345 3365 48385 3405
rect 50025 3365 50065 3405
rect 53300 3365 53340 3405
rect 54980 3365 55020 3405
rect 58255 3365 58295 3405
rect 59935 3365 59975 3405
rect 63210 3365 63250 3405
rect 64890 3365 64930 3405
rect 68165 3365 68205 3405
rect 69845 3365 69885 3405
rect 73120 3365 73160 3405
rect 74800 3365 74840 3405
rect 675 3080 715 3120
rect 675 2800 715 2835
rect 675 2450 715 2490
rect 1875 2800 1915 2835
rect 2355 2800 2395 2835
rect 3555 2800 3595 2835
rect 5630 3080 5670 3120
rect 5630 2800 5670 2835
rect 5630 2450 5670 2490
rect 6830 3080 6870 3120
rect 7310 3080 7350 3120
rect 6830 2800 6870 2835
rect 7310 2800 7350 2835
rect 6830 2450 6870 2490
rect 7310 2450 7350 2490
rect 8510 3080 8550 3120
rect 8510 2800 8550 2835
rect 8510 2450 8550 2490
rect 10585 3080 10625 3120
rect 10585 2800 10625 2835
rect 10585 2450 10625 2490
rect 11785 3080 11825 3120
rect 12265 3080 12305 3120
rect 11785 2800 11825 2835
rect 12265 2800 12305 2835
rect 11785 2450 11825 2490
rect 12265 2450 12305 2490
rect 13465 3080 13505 3120
rect 13465 2800 13505 2835
rect 13465 2450 13505 2490
rect 15540 3080 15580 3120
rect 15540 2800 15580 2835
rect 15540 2450 15580 2490
rect 16740 3080 16780 3120
rect 17220 3080 17260 3120
rect 16740 2800 16780 2835
rect 17220 2800 17260 2835
rect 16740 2450 16780 2490
rect 17220 2450 17260 2490
rect 18420 3080 18460 3120
rect 18420 2800 18460 2835
rect 18420 2450 18460 2490
rect 20495 3080 20535 3120
rect 20495 2800 20535 2835
rect 20495 2450 20535 2490
rect 21695 3080 21735 3120
rect 22175 3080 22215 3120
rect 21695 2800 21735 2835
rect 22175 2800 22215 2835
rect 21695 2450 21735 2490
rect 22175 2450 22215 2490
rect 23375 3080 23415 3120
rect 23375 2800 23415 2835
rect 23375 2450 23415 2490
rect 25450 3080 25490 3120
rect 25450 2800 25490 2835
rect 25450 2450 25490 2490
rect 26650 3080 26690 3120
rect 27130 3080 27170 3120
rect 26650 2800 26690 2835
rect 27130 2800 27170 2835
rect 26650 2450 26690 2490
rect 27130 2450 27170 2490
rect 28330 3080 28370 3120
rect 28330 2800 28370 2835
rect 28330 2450 28370 2490
rect 30405 3080 30445 3120
rect 30405 2800 30445 2835
rect 30405 2450 30445 2490
rect 31605 3080 31645 3120
rect 32085 3080 32125 3120
rect 31605 2800 31645 2835
rect 32085 2800 32125 2835
rect 31605 2450 31645 2490
rect 32085 2450 32125 2490
rect 33285 3080 33325 3120
rect 33285 2800 33325 2835
rect 33285 2450 33325 2490
rect 35360 3080 35400 3120
rect 35360 2800 35400 2835
rect 35360 2450 35400 2490
rect 36560 3080 36600 3120
rect 37040 3080 37080 3120
rect 36560 2800 36600 2835
rect 37040 2800 37080 2835
rect 36560 2450 36600 2490
rect 37040 2450 37080 2490
rect 38240 3080 38280 3120
rect 38240 2800 38280 2835
rect 38240 2450 38280 2490
rect 40315 3080 40355 3120
rect 40315 2800 40355 2835
rect 40315 2450 40355 2490
rect 41515 3080 41555 3120
rect 41995 3080 42035 3120
rect 41515 2800 41555 2835
rect 41995 2800 42035 2835
rect 41515 2450 41555 2490
rect 41995 2450 42035 2490
rect 43195 3080 43235 3120
rect 43195 2800 43235 2835
rect 43195 2450 43235 2490
rect 45270 3080 45310 3120
rect 45270 2800 45310 2835
rect 45270 2450 45310 2490
rect 46470 3080 46510 3120
rect 46950 3080 46990 3120
rect 46470 2800 46510 2835
rect 46950 2800 46990 2835
rect 46470 2450 46510 2490
rect 46950 2450 46990 2490
rect 48150 3080 48190 3120
rect 48150 2800 48190 2835
rect 48150 2450 48190 2490
rect 50225 3080 50265 3120
rect 50225 2800 50265 2835
rect 50225 2450 50265 2490
rect 51425 3080 51465 3120
rect 51905 3080 51945 3120
rect 51425 2800 51465 2835
rect 51905 2800 51945 2835
rect 51425 2450 51465 2490
rect 51905 2450 51945 2490
rect 53105 3080 53145 3120
rect 53105 2800 53145 2835
rect 53105 2450 53145 2490
rect 55180 3080 55220 3120
rect 55180 2800 55220 2835
rect 55180 2450 55220 2490
rect 56380 3080 56420 3120
rect 56860 3080 56900 3120
rect 56380 2800 56420 2835
rect 56860 2800 56900 2835
rect 56380 2450 56420 2490
rect 56860 2450 56900 2490
rect 58060 3080 58100 3120
rect 58060 2800 58100 2835
rect 58060 2450 58100 2490
rect 60135 3080 60175 3120
rect 60135 2800 60175 2835
rect 60135 2450 60175 2490
rect 61335 3080 61375 3120
rect 61815 3080 61855 3120
rect 61335 2800 61375 2835
rect 61815 2800 61855 2835
rect 61335 2450 61375 2490
rect 61815 2450 61855 2490
rect 63015 3080 63055 3120
rect 63015 2800 63055 2835
rect 63015 2450 63055 2490
rect 65090 3080 65130 3120
rect 65090 2800 65130 2835
rect 65090 2450 65130 2490
rect 66290 3080 66330 3120
rect 66770 3080 66810 3120
rect 66290 2800 66330 2835
rect 66770 2800 66810 2835
rect 66290 2450 66330 2490
rect 66770 2450 66810 2490
rect 67970 3080 68010 3120
rect 67970 2800 68010 2835
rect 67970 2450 68010 2490
rect 70045 3080 70085 3120
rect 70045 2800 70085 2835
rect 70045 2450 70085 2490
rect 71245 3080 71285 3120
rect 71725 3080 71765 3120
rect 71245 2800 71285 2835
rect 71725 2800 71765 2835
rect 71245 2450 71285 2490
rect 71725 2450 71765 2490
rect 72925 3080 72965 3120
rect 72925 2800 72965 2835
rect 72925 2450 72965 2490
rect 75000 3080 75040 3120
rect 75000 2800 75040 2835
rect 75000 2450 75040 2490
rect 76200 3080 76240 3120
rect 76680 3080 76720 3120
rect 76200 2800 76240 2835
rect 76680 2800 76720 2835
rect 76200 2450 76240 2490
rect 76680 2450 76720 2490
rect 77880 3080 77920 3120
rect 77880 2800 77920 2835
rect 77880 2450 77920 2490
rect 8705 2210 8745 2250
rect 10385 2210 10425 2250
rect 13660 2210 13700 2250
rect 15340 2210 15380 2250
rect 18615 2210 18655 2250
rect 20295 2210 20335 2250
rect 23570 2210 23610 2250
rect 25250 2210 25290 2250
rect 28525 2210 28565 2250
rect 30205 2210 30245 2250
rect 33480 2210 33520 2250
rect 35160 2210 35200 2250
rect 38435 2210 38475 2250
rect 40115 2210 40155 2250
rect 43390 2210 43430 2250
rect 45070 2210 45110 2250
rect 48345 2210 48385 2250
rect 50025 2210 50065 2250
rect 53300 2210 53340 2250
rect 54980 2210 55020 2250
rect 58255 2210 58295 2250
rect 59935 2210 59975 2250
rect 63210 2210 63250 2250
rect 64890 2210 64930 2250
rect 68165 2210 68205 2250
rect 69845 2210 69885 2250
rect 73120 2210 73160 2250
rect 74800 2210 74840 2250
rect 8705 290 8745 330
rect 10385 290 10425 330
rect 13660 290 13700 330
rect 15340 290 15380 330
rect 18615 290 18655 330
rect 20295 290 20335 330
rect 23570 290 23610 330
rect 25250 290 25290 330
rect 28525 290 28565 330
rect 30205 290 30245 330
rect 33480 290 33520 330
rect 35160 290 35200 330
rect 38435 290 38475 330
rect 40115 290 40155 330
rect 43390 290 43430 330
rect 45070 290 45110 330
rect 48345 290 48385 330
rect 50025 290 50065 330
rect 53300 290 53340 330
rect 54980 290 55020 330
rect 58255 290 58295 330
rect 59935 290 59975 330
rect 63210 290 63250 330
rect 64890 290 64930 330
rect 68165 290 68205 330
rect 69845 290 69885 330
rect 73120 290 73160 330
rect 74800 290 74840 330
<< metal1 >>
rect -345 12050 -185 12065
rect -345 11920 -330 12050
rect -200 11920 -185 12050
rect -345 11905 -185 11920
rect -345 11630 -280 11645
rect -345 11595 -330 11630
rect -295 11610 -280 11630
rect -295 11595 0 11610
rect -345 11580 0 11595
rect 4295 11580 4955 11610
rect 9250 11580 9910 11610
rect 14205 11580 14865 11610
rect 19160 11580 19820 11610
rect 24115 11580 24775 11610
rect 29070 11580 29730 11610
rect 34025 11580 34685 11610
rect 38980 11580 39640 11610
rect 43935 11580 44595 11610
rect 48890 11580 49550 11610
rect 53845 11580 54505 11610
rect 58800 11580 59460 11610
rect 63755 11580 64415 11610
rect 68710 11580 69370 11610
rect 73665 11580 74325 11610
rect 8690 11475 8775 11490
rect 8690 11435 8705 11475
rect 8745 11435 8775 11475
rect 8690 11420 8775 11435
rect 10355 11475 10440 11490
rect 10355 11435 10385 11475
rect 10425 11435 10440 11475
rect 10355 11420 10440 11435
rect 13645 11475 13730 11490
rect 13645 11435 13660 11475
rect 13700 11435 13730 11475
rect 13645 11420 13730 11435
rect 15310 11475 15395 11490
rect 15310 11435 15340 11475
rect 15380 11435 15395 11475
rect 15310 11420 15395 11435
rect 18600 11475 18685 11490
rect 18600 11435 18615 11475
rect 18655 11435 18685 11475
rect 18600 11420 18685 11435
rect 20265 11475 20350 11490
rect 20265 11435 20295 11475
rect 20335 11435 20350 11475
rect 20265 11420 20350 11435
rect 23555 11475 23640 11490
rect 23555 11435 23570 11475
rect 23610 11435 23640 11475
rect 23555 11420 23640 11435
rect 25220 11475 25305 11490
rect 25220 11435 25250 11475
rect 25290 11435 25305 11475
rect 25220 11420 25305 11435
rect 28510 11475 28595 11490
rect 28510 11435 28525 11475
rect 28565 11435 28595 11475
rect 28510 11420 28595 11435
rect 30175 11475 30260 11490
rect 30175 11435 30205 11475
rect 30245 11435 30260 11475
rect 30175 11420 30260 11435
rect 33465 11475 33550 11490
rect 33465 11435 33480 11475
rect 33520 11435 33550 11475
rect 33465 11420 33550 11435
rect 35130 11475 35215 11490
rect 35130 11435 35160 11475
rect 35200 11435 35215 11475
rect 35130 11420 35215 11435
rect 38420 11475 38505 11490
rect 38420 11435 38435 11475
rect 38475 11435 38505 11475
rect 38420 11420 38505 11435
rect 40085 11475 40170 11490
rect 40085 11435 40115 11475
rect 40155 11435 40170 11475
rect 40085 11420 40170 11435
rect 43375 11475 43460 11490
rect 43375 11435 43390 11475
rect 43430 11435 43460 11475
rect 43375 11420 43460 11435
rect 45040 11475 45125 11490
rect 45040 11435 45070 11475
rect 45110 11435 45125 11475
rect 45040 11420 45125 11435
rect 48330 11475 48415 11490
rect 48330 11435 48345 11475
rect 48385 11435 48415 11475
rect 48330 11420 48415 11435
rect 49995 11475 50080 11490
rect 49995 11435 50025 11475
rect 50065 11435 50080 11475
rect 49995 11420 50080 11435
rect 53285 11475 53370 11490
rect 53285 11435 53300 11475
rect 53340 11435 53370 11475
rect 53285 11420 53370 11435
rect 54950 11475 55035 11490
rect 54950 11435 54980 11475
rect 55020 11435 55035 11475
rect 54950 11420 55035 11435
rect 58240 11475 58325 11490
rect 58240 11435 58255 11475
rect 58295 11435 58325 11475
rect 58240 11420 58325 11435
rect 59905 11475 59990 11490
rect 59905 11435 59935 11475
rect 59975 11435 59990 11475
rect 59905 11420 59990 11435
rect 63195 11475 63280 11490
rect 63195 11435 63210 11475
rect 63250 11435 63280 11475
rect 63195 11420 63280 11435
rect 64860 11475 64945 11490
rect 64860 11435 64890 11475
rect 64930 11435 64945 11475
rect 64860 11420 64945 11435
rect 68150 11475 68235 11490
rect 68150 11435 68165 11475
rect 68205 11435 68235 11475
rect 68150 11420 68235 11435
rect 69815 11475 69900 11490
rect 69815 11435 69845 11475
rect 69885 11435 69900 11475
rect 69815 11420 69900 11435
rect 73105 11475 73190 11490
rect 73105 11435 73120 11475
rect 73160 11435 73190 11475
rect 73105 11420 73190 11435
rect 74770 11475 74855 11490
rect 74770 11435 74800 11475
rect 74840 11435 74855 11475
rect 74770 11420 74855 11435
rect 8690 9555 8775 9570
rect 8690 9515 8705 9555
rect 8745 9515 8775 9555
rect 8690 9500 8775 9515
rect 10355 9555 10440 9570
rect 10355 9515 10385 9555
rect 10425 9515 10440 9555
rect 10355 9500 10440 9515
rect 13645 9555 13730 9570
rect 13645 9515 13660 9555
rect 13700 9515 13730 9555
rect 13645 9500 13730 9515
rect 15310 9555 15395 9570
rect 15310 9515 15340 9555
rect 15380 9515 15395 9555
rect 15310 9500 15395 9515
rect 18600 9555 18685 9570
rect 18600 9515 18615 9555
rect 18655 9515 18685 9555
rect 18600 9500 18685 9515
rect 20265 9555 20350 9570
rect 20265 9515 20295 9555
rect 20335 9515 20350 9555
rect 20265 9500 20350 9515
rect 23555 9555 23640 9570
rect 23555 9515 23570 9555
rect 23610 9515 23640 9555
rect 23555 9500 23640 9515
rect 25220 9555 25305 9570
rect 25220 9515 25250 9555
rect 25290 9515 25305 9555
rect 25220 9500 25305 9515
rect 28510 9555 28595 9570
rect 28510 9515 28525 9555
rect 28565 9515 28595 9555
rect 28510 9500 28595 9515
rect 30175 9555 30260 9570
rect 30175 9515 30205 9555
rect 30245 9515 30260 9555
rect 30175 9500 30260 9515
rect 33465 9555 33550 9570
rect 33465 9515 33480 9555
rect 33520 9515 33550 9555
rect 33465 9500 33550 9515
rect 35130 9555 35215 9570
rect 35130 9515 35160 9555
rect 35200 9515 35215 9555
rect 35130 9500 35215 9515
rect 38420 9555 38505 9570
rect 38420 9515 38435 9555
rect 38475 9515 38505 9555
rect 38420 9500 38505 9515
rect 40085 9555 40170 9570
rect 40085 9515 40115 9555
rect 40155 9515 40170 9555
rect 40085 9500 40170 9515
rect 43375 9555 43460 9570
rect 43375 9515 43390 9555
rect 43430 9515 43460 9555
rect 43375 9500 43460 9515
rect 45040 9555 45125 9570
rect 45040 9515 45070 9555
rect 45110 9515 45125 9555
rect 45040 9500 45125 9515
rect 48330 9555 48415 9570
rect 48330 9515 48345 9555
rect 48385 9515 48415 9555
rect 48330 9500 48415 9515
rect 49995 9555 50080 9570
rect 49995 9515 50025 9555
rect 50065 9515 50080 9555
rect 49995 9500 50080 9515
rect 53285 9555 53370 9570
rect 53285 9515 53300 9555
rect 53340 9515 53370 9555
rect 53285 9500 53370 9515
rect 54950 9555 55035 9570
rect 54950 9515 54980 9555
rect 55020 9515 55035 9555
rect 54950 9500 55035 9515
rect 58240 9555 58325 9570
rect 58240 9515 58255 9555
rect 58295 9515 58325 9555
rect 58240 9500 58325 9515
rect 59905 9555 59990 9570
rect 59905 9515 59935 9555
rect 59975 9515 59990 9555
rect 59905 9500 59990 9515
rect 63195 9555 63280 9570
rect 63195 9515 63210 9555
rect 63250 9515 63280 9555
rect 63195 9500 63280 9515
rect 64860 9555 64945 9570
rect 64860 9515 64890 9555
rect 64930 9515 64945 9555
rect 64860 9500 64945 9515
rect 68150 9555 68235 9570
rect 68150 9515 68165 9555
rect 68205 9515 68235 9555
rect 68150 9500 68235 9515
rect 69815 9555 69900 9570
rect 69815 9515 69845 9555
rect 69885 9515 69900 9555
rect 69815 9500 69900 9515
rect 73105 9555 73190 9570
rect 73105 9515 73120 9555
rect 73160 9515 73190 9555
rect 73105 9500 73190 9515
rect 74770 9555 74855 9570
rect 74770 9515 74800 9555
rect 74840 9515 74855 9555
rect 74770 9500 74855 9515
rect 15 9410 80 9425
rect 15 9375 30 9410
rect 65 9375 80 9410
rect 15 9360 80 9375
rect 4365 9360 4970 9390
rect 9320 9360 9925 9390
rect 14275 9360 14880 9390
rect 19230 9360 19835 9390
rect 24185 9360 24790 9390
rect 29140 9360 29745 9390
rect 34095 9360 34700 9390
rect 39050 9360 39655 9390
rect 44005 9360 44610 9390
rect 48960 9360 49565 9390
rect 53915 9360 54520 9390
rect 58870 9360 59475 9390
rect 63825 9360 64430 9390
rect 68780 9360 69385 9390
rect 73735 9360 74340 9390
rect 5615 9270 5685 9285
rect 5615 9230 5630 9270
rect 5670 9230 5685 9270
rect 5615 9200 5685 9230
rect 6815 9270 6885 9285
rect 6815 9230 6830 9270
rect 6870 9230 6885 9270
rect 6815 9200 6885 9230
rect 7295 9270 7365 9285
rect 7295 9230 7310 9270
rect 7350 9230 7365 9270
rect 7295 9200 7365 9230
rect 8495 9270 8565 9285
rect 8495 9230 8510 9270
rect 8550 9230 8565 9270
rect 8495 9200 8565 9230
rect 10570 9270 10640 9285
rect 10570 9230 10585 9270
rect 10625 9230 10640 9270
rect 10570 9200 10640 9230
rect 11770 9270 11840 9285
rect 11770 9230 11785 9270
rect 11825 9230 11840 9270
rect 11770 9200 11840 9230
rect 12250 9270 12320 9285
rect 12250 9230 12265 9270
rect 12305 9230 12320 9270
rect 12250 9200 12320 9230
rect 13450 9270 13520 9285
rect 13450 9230 13465 9270
rect 13505 9230 13520 9270
rect 13450 9200 13520 9230
rect 15525 9270 15595 9285
rect 15525 9230 15540 9270
rect 15580 9230 15595 9270
rect 15525 9200 15595 9230
rect 16725 9270 16795 9285
rect 16725 9230 16740 9270
rect 16780 9230 16795 9270
rect 16725 9200 16795 9230
rect 17205 9270 17275 9285
rect 17205 9230 17220 9270
rect 17260 9230 17275 9270
rect 17205 9200 17275 9230
rect 18405 9270 18475 9285
rect 18405 9230 18420 9270
rect 18460 9230 18475 9270
rect 18405 9200 18475 9230
rect 20480 9270 20550 9285
rect 20480 9230 20495 9270
rect 20535 9230 20550 9270
rect 20480 9200 20550 9230
rect 21680 9270 21750 9285
rect 21680 9230 21695 9270
rect 21735 9230 21750 9270
rect 21680 9200 21750 9230
rect 22160 9270 22230 9285
rect 22160 9230 22175 9270
rect 22215 9230 22230 9270
rect 22160 9200 22230 9230
rect 23360 9270 23430 9285
rect 23360 9230 23375 9270
rect 23415 9230 23430 9270
rect 23360 9200 23430 9230
rect 25435 9270 25505 9285
rect 25435 9230 25450 9270
rect 25490 9230 25505 9270
rect 25435 9200 25505 9230
rect 26635 9270 26705 9285
rect 26635 9230 26650 9270
rect 26690 9230 26705 9270
rect 26635 9200 26705 9230
rect 27115 9270 27185 9285
rect 27115 9230 27130 9270
rect 27170 9230 27185 9270
rect 27115 9200 27185 9230
rect 28315 9270 28385 9285
rect 28315 9230 28330 9270
rect 28370 9230 28385 9270
rect 28315 9200 28385 9230
rect 30390 9270 30460 9285
rect 30390 9230 30405 9270
rect 30445 9230 30460 9270
rect 30390 9200 30460 9230
rect 31590 9270 31660 9285
rect 31590 9230 31605 9270
rect 31645 9230 31660 9270
rect 31590 9200 31660 9230
rect 32070 9270 32140 9285
rect 32070 9230 32085 9270
rect 32125 9230 32140 9270
rect 32070 9200 32140 9230
rect 33270 9270 33340 9285
rect 33270 9230 33285 9270
rect 33325 9230 33340 9270
rect 33270 9200 33340 9230
rect 35345 9270 35415 9285
rect 35345 9230 35360 9270
rect 35400 9230 35415 9270
rect 35345 9200 35415 9230
rect 36545 9270 36615 9285
rect 36545 9230 36560 9270
rect 36600 9230 36615 9270
rect 36545 9200 36615 9230
rect 37025 9270 37095 9285
rect 37025 9230 37040 9270
rect 37080 9230 37095 9270
rect 37025 9200 37095 9230
rect 38225 9270 38295 9285
rect 38225 9230 38240 9270
rect 38280 9230 38295 9270
rect 38225 9200 38295 9230
rect 40300 9270 40370 9285
rect 40300 9230 40315 9270
rect 40355 9230 40370 9270
rect 40300 9200 40370 9230
rect 41500 9270 41570 9285
rect 41500 9230 41515 9270
rect 41555 9230 41570 9270
rect 41500 9200 41570 9230
rect 41980 9270 42050 9285
rect 41980 9230 41995 9270
rect 42035 9230 42050 9270
rect 41980 9200 42050 9230
rect 43180 9270 43250 9285
rect 43180 9230 43195 9270
rect 43235 9230 43250 9270
rect 43180 9200 43250 9230
rect 45255 9270 45325 9285
rect 45255 9230 45270 9270
rect 45310 9230 45325 9270
rect 45255 9200 45325 9230
rect 46455 9270 46525 9285
rect 46455 9230 46470 9270
rect 46510 9230 46525 9270
rect 46455 9200 46525 9230
rect 46935 9270 47005 9285
rect 46935 9230 46950 9270
rect 46990 9230 47005 9270
rect 46935 9200 47005 9230
rect 48135 9270 48205 9285
rect 48135 9230 48150 9270
rect 48190 9230 48205 9270
rect 48135 9200 48205 9230
rect 50210 9270 50280 9285
rect 50210 9230 50225 9270
rect 50265 9230 50280 9270
rect 50210 9200 50280 9230
rect 51410 9270 51480 9285
rect 51410 9230 51425 9270
rect 51465 9230 51480 9270
rect 51410 9200 51480 9230
rect 51890 9270 51960 9285
rect 51890 9230 51905 9270
rect 51945 9230 51960 9270
rect 51890 9200 51960 9230
rect 53090 9270 53160 9285
rect 53090 9230 53105 9270
rect 53145 9230 53160 9270
rect 53090 9200 53160 9230
rect 55165 9270 55235 9285
rect 55165 9230 55180 9270
rect 55220 9230 55235 9270
rect 55165 9200 55235 9230
rect 56365 9270 56435 9285
rect 56365 9230 56380 9270
rect 56420 9230 56435 9270
rect 56365 9200 56435 9230
rect 56845 9270 56915 9285
rect 56845 9230 56860 9270
rect 56900 9230 56915 9270
rect 56845 9200 56915 9230
rect 58045 9270 58115 9285
rect 58045 9230 58060 9270
rect 58100 9230 58115 9270
rect 58045 9200 58115 9230
rect 60120 9270 60190 9285
rect 60120 9230 60135 9270
rect 60175 9230 60190 9270
rect 60120 9200 60190 9230
rect 61320 9270 61390 9285
rect 61320 9230 61335 9270
rect 61375 9230 61390 9270
rect 61320 9200 61390 9230
rect 61800 9270 61870 9285
rect 61800 9230 61815 9270
rect 61855 9230 61870 9270
rect 61800 9200 61870 9230
rect 63000 9270 63070 9285
rect 63000 9230 63015 9270
rect 63055 9230 63070 9270
rect 63000 9200 63070 9230
rect 65075 9270 65145 9285
rect 65075 9230 65090 9270
rect 65130 9230 65145 9270
rect 65075 9200 65145 9230
rect 66275 9270 66345 9285
rect 66275 9230 66290 9270
rect 66330 9230 66345 9270
rect 66275 9200 66345 9230
rect 66755 9270 66825 9285
rect 66755 9230 66770 9270
rect 66810 9230 66825 9270
rect 66755 9200 66825 9230
rect 67955 9270 68025 9285
rect 67955 9230 67970 9270
rect 68010 9230 68025 9270
rect 67955 9200 68025 9230
rect 70030 9270 70100 9285
rect 70030 9230 70045 9270
rect 70085 9230 70100 9270
rect 70030 9200 70100 9230
rect 71230 9270 71300 9285
rect 71230 9230 71245 9270
rect 71285 9230 71300 9270
rect 71230 9200 71300 9230
rect 71710 9270 71780 9285
rect 71710 9230 71725 9270
rect 71765 9230 71780 9270
rect 71710 9200 71780 9230
rect 72910 9270 72980 9285
rect 72910 9230 72925 9270
rect 72965 9230 72980 9270
rect 72910 9200 72980 9230
rect 74985 9270 75055 9285
rect 74985 9230 75000 9270
rect 75040 9230 75055 9270
rect 74985 9200 75055 9230
rect 76185 9270 76255 9285
rect 76185 9230 76200 9270
rect 76240 9230 76255 9270
rect 76185 9200 76255 9230
rect 76665 9270 76735 9285
rect 76665 9230 76680 9270
rect 76720 9230 76735 9270
rect 76665 9200 76735 9230
rect 77865 9270 77935 9285
rect 77865 9230 77880 9270
rect 77920 9230 77935 9270
rect 77865 9200 77935 9230
rect 660 8935 77935 8950
rect 660 8900 675 8935
rect 715 8900 1875 8935
rect 1915 8900 2355 8935
rect 2395 8900 3555 8935
rect 3595 8900 5630 8935
rect 5670 8900 6830 8935
rect 6870 8900 7310 8935
rect 7350 8900 8510 8935
rect 8550 8900 10585 8935
rect 10625 8900 11785 8935
rect 11825 8900 12265 8935
rect 12305 8900 13465 8935
rect 13505 8900 15540 8935
rect 15580 8900 16740 8935
rect 16780 8900 17220 8935
rect 17260 8900 18420 8935
rect 18460 8900 20495 8935
rect 20535 8900 21695 8935
rect 21735 8900 22175 8935
rect 22215 8900 23375 8935
rect 23415 8900 25450 8935
rect 25490 8900 26650 8935
rect 26690 8900 27130 8935
rect 27170 8900 28330 8935
rect 28370 8900 30405 8935
rect 30445 8900 31605 8935
rect 31645 8900 32085 8935
rect 32125 8900 33285 8935
rect 33325 8900 35360 8935
rect 35400 8900 36560 8935
rect 36600 8900 37040 8935
rect 37080 8900 38240 8935
rect 38280 8900 40315 8935
rect 40355 8900 41515 8935
rect 41555 8900 41995 8935
rect 42035 8900 43195 8935
rect 43235 8900 45270 8935
rect 45310 8900 46470 8935
rect 46510 8900 46950 8935
rect 46990 8900 48150 8935
rect 48190 8900 50225 8935
rect 50265 8900 51425 8935
rect 51465 8900 51905 8935
rect 51945 8900 53105 8935
rect 53145 8900 55180 8935
rect 55220 8900 56380 8935
rect 56420 8900 56860 8935
rect 56900 8900 58060 8935
rect 58100 8900 60135 8935
rect 60175 8900 61335 8935
rect 61375 8900 61815 8935
rect 61855 8900 63015 8935
rect 63055 8900 65090 8935
rect 65130 8900 66290 8935
rect 66330 8900 66770 8935
rect 66810 8900 67970 8935
rect 68010 8900 70045 8935
rect 70085 8900 71245 8935
rect 71285 8900 71725 8935
rect 71765 8900 72925 8935
rect 72965 8900 75000 8935
rect 75040 8900 76200 8935
rect 76240 8900 76680 8935
rect 76720 8900 77880 8935
rect 77920 8900 77935 8935
rect 660 8885 77935 8900
rect 5615 8640 5685 8670
rect 5615 8600 5630 8640
rect 5670 8600 5685 8640
rect 5615 8585 5685 8600
rect 6815 8640 6885 8670
rect 6815 8600 6830 8640
rect 6870 8600 6885 8640
rect 6815 8585 6885 8600
rect 7295 8640 7365 8670
rect 7295 8600 7310 8640
rect 7350 8600 7365 8640
rect 7295 8585 7365 8600
rect 8495 8640 8565 8670
rect 8495 8600 8510 8640
rect 8550 8600 8565 8640
rect 8495 8585 8565 8600
rect 10570 8640 10640 8670
rect 10570 8600 10585 8640
rect 10625 8600 10640 8640
rect 10570 8585 10640 8600
rect 11770 8640 11840 8670
rect 11770 8600 11785 8640
rect 11825 8600 11840 8640
rect 11770 8585 11840 8600
rect 12250 8640 12320 8670
rect 12250 8600 12265 8640
rect 12305 8600 12320 8640
rect 12250 8585 12320 8600
rect 13450 8640 13520 8670
rect 13450 8600 13465 8640
rect 13505 8600 13520 8640
rect 13450 8585 13520 8600
rect 15525 8640 15595 8670
rect 15525 8600 15540 8640
rect 15580 8600 15595 8640
rect 15525 8585 15595 8600
rect 16725 8640 16795 8670
rect 16725 8600 16740 8640
rect 16780 8600 16795 8640
rect 16725 8585 16795 8600
rect 17205 8640 17275 8670
rect 17205 8600 17220 8640
rect 17260 8600 17275 8640
rect 17205 8585 17275 8600
rect 18405 8640 18475 8670
rect 18405 8600 18420 8640
rect 18460 8600 18475 8640
rect 18405 8585 18475 8600
rect 20480 8640 20550 8670
rect 20480 8600 20495 8640
rect 20535 8600 20550 8640
rect 20480 8585 20550 8600
rect 21680 8640 21750 8670
rect 21680 8600 21695 8640
rect 21735 8600 21750 8640
rect 21680 8585 21750 8600
rect 22160 8640 22230 8670
rect 22160 8600 22175 8640
rect 22215 8600 22230 8640
rect 22160 8585 22230 8600
rect 23360 8640 23430 8670
rect 23360 8600 23375 8640
rect 23415 8600 23430 8640
rect 23360 8585 23430 8600
rect 25435 8640 25505 8670
rect 25435 8600 25450 8640
rect 25490 8600 25505 8640
rect 25435 8585 25505 8600
rect 26635 8640 26705 8670
rect 26635 8600 26650 8640
rect 26690 8600 26705 8640
rect 26635 8585 26705 8600
rect 27115 8640 27185 8670
rect 27115 8600 27130 8640
rect 27170 8600 27185 8640
rect 27115 8585 27185 8600
rect 28315 8640 28385 8670
rect 28315 8600 28330 8640
rect 28370 8600 28385 8640
rect 28315 8585 28385 8600
rect 30390 8640 30460 8670
rect 30390 8600 30405 8640
rect 30445 8600 30460 8640
rect 30390 8585 30460 8600
rect 31590 8640 31660 8670
rect 31590 8600 31605 8640
rect 31645 8600 31660 8640
rect 31590 8585 31660 8600
rect 32070 8640 32140 8670
rect 32070 8600 32085 8640
rect 32125 8600 32140 8640
rect 32070 8585 32140 8600
rect 33270 8640 33340 8670
rect 33270 8600 33285 8640
rect 33325 8600 33340 8640
rect 33270 8585 33340 8600
rect 35345 8640 35415 8670
rect 35345 8600 35360 8640
rect 35400 8600 35415 8640
rect 35345 8585 35415 8600
rect 36545 8640 36615 8670
rect 36545 8600 36560 8640
rect 36600 8600 36615 8640
rect 36545 8585 36615 8600
rect 37025 8640 37095 8670
rect 37025 8600 37040 8640
rect 37080 8600 37095 8640
rect 37025 8585 37095 8600
rect 38225 8640 38295 8670
rect 38225 8600 38240 8640
rect 38280 8600 38295 8640
rect 38225 8585 38295 8600
rect 40300 8640 40370 8670
rect 40300 8600 40315 8640
rect 40355 8600 40370 8640
rect 40300 8585 40370 8600
rect 41500 8640 41570 8670
rect 41500 8600 41515 8640
rect 41555 8600 41570 8640
rect 41500 8585 41570 8600
rect 41980 8640 42050 8670
rect 41980 8600 41995 8640
rect 42035 8600 42050 8640
rect 41980 8585 42050 8600
rect 43180 8640 43250 8670
rect 43180 8600 43195 8640
rect 43235 8600 43250 8640
rect 43180 8585 43250 8600
rect 45255 8640 45325 8670
rect 45255 8600 45270 8640
rect 45310 8600 45325 8640
rect 45255 8585 45325 8600
rect 46455 8640 46525 8670
rect 46455 8600 46470 8640
rect 46510 8600 46525 8640
rect 46455 8585 46525 8600
rect 46935 8640 47005 8670
rect 46935 8600 46950 8640
rect 46990 8600 47005 8640
rect 46935 8585 47005 8600
rect 48135 8640 48205 8670
rect 48135 8600 48150 8640
rect 48190 8600 48205 8640
rect 48135 8585 48205 8600
rect 50210 8640 50280 8670
rect 50210 8600 50225 8640
rect 50265 8600 50280 8640
rect 50210 8585 50280 8600
rect 51410 8640 51480 8670
rect 51410 8600 51425 8640
rect 51465 8600 51480 8640
rect 51410 8585 51480 8600
rect 51890 8640 51960 8670
rect 51890 8600 51905 8640
rect 51945 8600 51960 8640
rect 51890 8585 51960 8600
rect 53090 8640 53160 8670
rect 53090 8600 53105 8640
rect 53145 8600 53160 8640
rect 53090 8585 53160 8600
rect 55165 8640 55235 8670
rect 55165 8600 55180 8640
rect 55220 8600 55235 8640
rect 55165 8585 55235 8600
rect 56365 8640 56435 8670
rect 56365 8600 56380 8640
rect 56420 8600 56435 8640
rect 56365 8585 56435 8600
rect 56845 8640 56915 8670
rect 56845 8600 56860 8640
rect 56900 8600 56915 8640
rect 56845 8585 56915 8600
rect 58045 8640 58115 8670
rect 58045 8600 58060 8640
rect 58100 8600 58115 8640
rect 58045 8585 58115 8600
rect 60120 8640 60190 8670
rect 60120 8600 60135 8640
rect 60175 8600 60190 8640
rect 60120 8585 60190 8600
rect 61320 8640 61390 8670
rect 61320 8600 61335 8640
rect 61375 8600 61390 8640
rect 61320 8585 61390 8600
rect 61800 8640 61870 8670
rect 61800 8600 61815 8640
rect 61855 8600 61870 8640
rect 61800 8585 61870 8600
rect 63000 8640 63070 8670
rect 63000 8600 63015 8640
rect 63055 8600 63070 8640
rect 63000 8585 63070 8600
rect 65075 8640 65145 8670
rect 65075 8600 65090 8640
rect 65130 8600 65145 8640
rect 65075 8585 65145 8600
rect 66275 8640 66345 8670
rect 66275 8600 66290 8640
rect 66330 8600 66345 8640
rect 66275 8585 66345 8600
rect 66755 8640 66825 8670
rect 66755 8600 66770 8640
rect 66810 8600 66825 8640
rect 66755 8585 66825 8600
rect 67955 8640 68025 8670
rect 67955 8600 67970 8640
rect 68010 8600 68025 8640
rect 67955 8585 68025 8600
rect 70030 8640 70100 8670
rect 70030 8600 70045 8640
rect 70085 8600 70100 8640
rect 70030 8585 70100 8600
rect 71230 8640 71300 8670
rect 71230 8600 71245 8640
rect 71285 8600 71300 8640
rect 71230 8585 71300 8600
rect 71710 8640 71780 8670
rect 71710 8600 71725 8640
rect 71765 8600 71780 8640
rect 71710 8585 71780 8600
rect 72910 8640 72980 8670
rect 72910 8600 72925 8640
rect 72965 8600 72980 8640
rect 72910 8585 72980 8600
rect 74985 8640 75055 8670
rect 74985 8600 75000 8640
rect 75040 8600 75055 8640
rect 74985 8585 75055 8600
rect 76185 8640 76255 8670
rect 76185 8600 76200 8640
rect 76240 8600 76255 8640
rect 76185 8585 76255 8600
rect 76665 8640 76735 8670
rect 76665 8600 76680 8640
rect 76720 8600 76735 8640
rect 76665 8585 76735 8600
rect 77865 8640 77935 8670
rect 77865 8600 77880 8640
rect 77920 8600 77935 8640
rect 77865 8585 77935 8600
rect -345 8555 -280 8570
rect -345 8520 -330 8555
rect -295 8535 -280 8555
rect -295 8520 0 8535
rect -345 8505 0 8520
rect 4295 8505 4955 8535
rect 9250 8505 9910 8535
rect 14205 8505 14865 8535
rect 19160 8505 19820 8535
rect 24115 8505 24775 8535
rect 29070 8505 29730 8535
rect 34025 8505 34685 8535
rect 38980 8505 39640 8535
rect 43935 8505 44595 8535
rect 48890 8505 49550 8535
rect 53845 8505 54505 8535
rect 58800 8505 59460 8535
rect 63755 8505 64415 8535
rect 68710 8505 69370 8535
rect 73665 8505 74325 8535
rect 8690 8400 8775 8415
rect 8690 8360 8705 8400
rect 8745 8360 8775 8400
rect 8690 8345 8775 8360
rect 10355 8400 10440 8415
rect 10355 8360 10385 8400
rect 10425 8360 10440 8400
rect 10355 8345 10440 8360
rect 13645 8400 13730 8415
rect 13645 8360 13660 8400
rect 13700 8360 13730 8400
rect 13645 8345 13730 8360
rect 15310 8400 15395 8415
rect 15310 8360 15340 8400
rect 15380 8360 15395 8400
rect 15310 8345 15395 8360
rect 18600 8400 18685 8415
rect 18600 8360 18615 8400
rect 18655 8360 18685 8400
rect 18600 8345 18685 8360
rect 20265 8400 20350 8415
rect 20265 8360 20295 8400
rect 20335 8360 20350 8400
rect 20265 8345 20350 8360
rect 23555 8400 23640 8415
rect 23555 8360 23570 8400
rect 23610 8360 23640 8400
rect 23555 8345 23640 8360
rect 25220 8400 25305 8415
rect 25220 8360 25250 8400
rect 25290 8360 25305 8400
rect 25220 8345 25305 8360
rect 28510 8400 28595 8415
rect 28510 8360 28525 8400
rect 28565 8360 28595 8400
rect 28510 8345 28595 8360
rect 30175 8400 30260 8415
rect 30175 8360 30205 8400
rect 30245 8360 30260 8400
rect 30175 8345 30260 8360
rect 33465 8400 33550 8415
rect 33465 8360 33480 8400
rect 33520 8360 33550 8400
rect 33465 8345 33550 8360
rect 35130 8400 35215 8415
rect 35130 8360 35160 8400
rect 35200 8360 35215 8400
rect 35130 8345 35215 8360
rect 38420 8400 38505 8415
rect 38420 8360 38435 8400
rect 38475 8360 38505 8400
rect 38420 8345 38505 8360
rect 40085 8400 40170 8415
rect 40085 8360 40115 8400
rect 40155 8360 40170 8400
rect 40085 8345 40170 8360
rect 43375 8400 43460 8415
rect 43375 8360 43390 8400
rect 43430 8360 43460 8400
rect 43375 8345 43460 8360
rect 45040 8400 45125 8415
rect 45040 8360 45070 8400
rect 45110 8360 45125 8400
rect 45040 8345 45125 8360
rect 48330 8400 48415 8415
rect 48330 8360 48345 8400
rect 48385 8360 48415 8400
rect 48330 8345 48415 8360
rect 49995 8400 50080 8415
rect 49995 8360 50025 8400
rect 50065 8360 50080 8400
rect 49995 8345 50080 8360
rect 53285 8400 53370 8415
rect 53285 8360 53300 8400
rect 53340 8360 53370 8400
rect 53285 8345 53370 8360
rect 54950 8400 55035 8415
rect 54950 8360 54980 8400
rect 55020 8360 55035 8400
rect 54950 8345 55035 8360
rect 58240 8400 58325 8415
rect 58240 8360 58255 8400
rect 58295 8360 58325 8400
rect 58240 8345 58325 8360
rect 59905 8400 59990 8415
rect 59905 8360 59935 8400
rect 59975 8360 59990 8400
rect 59905 8345 59990 8360
rect 63195 8400 63280 8415
rect 63195 8360 63210 8400
rect 63250 8360 63280 8400
rect 63195 8345 63280 8360
rect 64860 8400 64945 8415
rect 64860 8360 64890 8400
rect 64930 8360 64945 8400
rect 64860 8345 64945 8360
rect 68150 8400 68235 8415
rect 68150 8360 68165 8400
rect 68205 8360 68235 8400
rect 68150 8345 68235 8360
rect 69815 8400 69900 8415
rect 69815 8360 69845 8400
rect 69885 8360 69900 8400
rect 69815 8345 69900 8360
rect 73105 8400 73190 8415
rect 73105 8360 73120 8400
rect 73160 8360 73190 8400
rect 73105 8345 73190 8360
rect 74770 8400 74855 8415
rect 74770 8360 74800 8400
rect 74840 8360 74855 8400
rect 74770 8345 74855 8360
rect 8690 6480 8775 6495
rect 8690 6440 8705 6480
rect 8745 6440 8775 6480
rect 8690 6425 8775 6440
rect 10355 6480 10440 6495
rect 10355 6440 10385 6480
rect 10425 6440 10440 6480
rect 10355 6425 10440 6440
rect 13645 6480 13730 6495
rect 13645 6440 13660 6480
rect 13700 6440 13730 6480
rect 13645 6425 13730 6440
rect 15310 6480 15395 6495
rect 15310 6440 15340 6480
rect 15380 6440 15395 6480
rect 15310 6425 15395 6440
rect 18600 6480 18685 6495
rect 18600 6440 18615 6480
rect 18655 6440 18685 6480
rect 18600 6425 18685 6440
rect 20265 6480 20350 6495
rect 20265 6440 20295 6480
rect 20335 6440 20350 6480
rect 20265 6425 20350 6440
rect 23555 6480 23640 6495
rect 23555 6440 23570 6480
rect 23610 6440 23640 6480
rect 23555 6425 23640 6440
rect 25220 6480 25305 6495
rect 25220 6440 25250 6480
rect 25290 6440 25305 6480
rect 25220 6425 25305 6440
rect 28510 6480 28595 6495
rect 28510 6440 28525 6480
rect 28565 6440 28595 6480
rect 28510 6425 28595 6440
rect 30175 6480 30260 6495
rect 30175 6440 30205 6480
rect 30245 6440 30260 6480
rect 30175 6425 30260 6440
rect 33465 6480 33550 6495
rect 33465 6440 33480 6480
rect 33520 6440 33550 6480
rect 33465 6425 33550 6440
rect 35130 6480 35215 6495
rect 35130 6440 35160 6480
rect 35200 6440 35215 6480
rect 35130 6425 35215 6440
rect 38420 6480 38505 6495
rect 38420 6440 38435 6480
rect 38475 6440 38505 6480
rect 38420 6425 38505 6440
rect 40085 6480 40170 6495
rect 40085 6440 40115 6480
rect 40155 6440 40170 6480
rect 40085 6425 40170 6440
rect 43375 6480 43460 6495
rect 43375 6440 43390 6480
rect 43430 6440 43460 6480
rect 43375 6425 43460 6440
rect 45040 6480 45125 6495
rect 45040 6440 45070 6480
rect 45110 6440 45125 6480
rect 45040 6425 45125 6440
rect 48330 6480 48415 6495
rect 48330 6440 48345 6480
rect 48385 6440 48415 6480
rect 48330 6425 48415 6440
rect 49995 6480 50080 6495
rect 49995 6440 50025 6480
rect 50065 6440 50080 6480
rect 49995 6425 50080 6440
rect 53285 6480 53370 6495
rect 53285 6440 53300 6480
rect 53340 6440 53370 6480
rect 53285 6425 53370 6440
rect 54950 6480 55035 6495
rect 54950 6440 54980 6480
rect 55020 6440 55035 6480
rect 54950 6425 55035 6440
rect 58240 6480 58325 6495
rect 58240 6440 58255 6480
rect 58295 6440 58325 6480
rect 58240 6425 58325 6440
rect 59905 6480 59990 6495
rect 59905 6440 59935 6480
rect 59975 6440 59990 6480
rect 59905 6425 59990 6440
rect 63195 6480 63280 6495
rect 63195 6440 63210 6480
rect 63250 6440 63280 6480
rect 63195 6425 63280 6440
rect 64860 6480 64945 6495
rect 64860 6440 64890 6480
rect 64930 6440 64945 6480
rect 64860 6425 64945 6440
rect 68150 6480 68235 6495
rect 68150 6440 68165 6480
rect 68205 6440 68235 6480
rect 68150 6425 68235 6440
rect 69815 6480 69900 6495
rect 69815 6440 69845 6480
rect 69885 6440 69900 6480
rect 69815 6425 69900 6440
rect 73105 6480 73190 6495
rect 73105 6440 73120 6480
rect 73160 6440 73190 6480
rect 73105 6425 73190 6440
rect 74770 6480 74855 6495
rect 74770 6440 74800 6480
rect 74840 6440 74855 6480
rect 74770 6425 74855 6440
rect 15 6335 80 6350
rect 15 6300 30 6335
rect 65 6300 80 6335
rect 15 6285 80 6300
rect 4365 6285 4970 6315
rect 9320 6285 9925 6315
rect 14275 6285 14880 6315
rect 19230 6285 19835 6315
rect 24185 6285 24790 6315
rect 29140 6285 29745 6315
rect 34095 6285 34700 6315
rect 39050 6285 39655 6315
rect 44005 6285 44610 6315
rect 48960 6285 49565 6315
rect 53915 6285 54520 6315
rect 58870 6285 59475 6315
rect 63825 6285 64430 6315
rect 68780 6285 69385 6315
rect 73735 6285 74340 6315
rect 5615 6195 5685 6210
rect 5615 6155 5630 6195
rect 5670 6155 5685 6195
rect 5615 6125 5685 6155
rect 6815 6195 6885 6210
rect 6815 6155 6830 6195
rect 6870 6155 6885 6195
rect 6815 6125 6885 6155
rect 7295 6195 7365 6210
rect 7295 6155 7310 6195
rect 7350 6155 7365 6195
rect 7295 6125 7365 6155
rect 8495 6195 8565 6210
rect 8495 6155 8510 6195
rect 8550 6155 8565 6195
rect 8495 6125 8565 6155
rect 10570 6195 10640 6210
rect 10570 6155 10585 6195
rect 10625 6155 10640 6195
rect 10570 6125 10640 6155
rect 11770 6195 11840 6210
rect 11770 6155 11785 6195
rect 11825 6155 11840 6195
rect 11770 6125 11840 6155
rect 12250 6195 12320 6210
rect 12250 6155 12265 6195
rect 12305 6155 12320 6195
rect 12250 6125 12320 6155
rect 13450 6195 13520 6210
rect 13450 6155 13465 6195
rect 13505 6155 13520 6195
rect 13450 6125 13520 6155
rect 15525 6195 15595 6210
rect 15525 6155 15540 6195
rect 15580 6155 15595 6195
rect 15525 6125 15595 6155
rect 16725 6195 16795 6210
rect 16725 6155 16740 6195
rect 16780 6155 16795 6195
rect 16725 6125 16795 6155
rect 17205 6195 17275 6210
rect 17205 6155 17220 6195
rect 17260 6155 17275 6195
rect 17205 6125 17275 6155
rect 18405 6195 18475 6210
rect 18405 6155 18420 6195
rect 18460 6155 18475 6195
rect 18405 6125 18475 6155
rect 20480 6195 20550 6210
rect 20480 6155 20495 6195
rect 20535 6155 20550 6195
rect 20480 6125 20550 6155
rect 21680 6195 21750 6210
rect 21680 6155 21695 6195
rect 21735 6155 21750 6195
rect 21680 6125 21750 6155
rect 22160 6195 22230 6210
rect 22160 6155 22175 6195
rect 22215 6155 22230 6195
rect 22160 6125 22230 6155
rect 23360 6195 23430 6210
rect 23360 6155 23375 6195
rect 23415 6155 23430 6195
rect 23360 6125 23430 6155
rect 25435 6195 25505 6210
rect 25435 6155 25450 6195
rect 25490 6155 25505 6195
rect 25435 6125 25505 6155
rect 26635 6195 26705 6210
rect 26635 6155 26650 6195
rect 26690 6155 26705 6195
rect 26635 6125 26705 6155
rect 27115 6195 27185 6210
rect 27115 6155 27130 6195
rect 27170 6155 27185 6195
rect 27115 6125 27185 6155
rect 28315 6195 28385 6210
rect 28315 6155 28330 6195
rect 28370 6155 28385 6195
rect 28315 6125 28385 6155
rect 30390 6195 30460 6210
rect 30390 6155 30405 6195
rect 30445 6155 30460 6195
rect 30390 6125 30460 6155
rect 31590 6195 31660 6210
rect 31590 6155 31605 6195
rect 31645 6155 31660 6195
rect 31590 6125 31660 6155
rect 32070 6195 32140 6210
rect 32070 6155 32085 6195
rect 32125 6155 32140 6195
rect 32070 6125 32140 6155
rect 33270 6195 33340 6210
rect 33270 6155 33285 6195
rect 33325 6155 33340 6195
rect 33270 6125 33340 6155
rect 35345 6195 35415 6210
rect 35345 6155 35360 6195
rect 35400 6155 35415 6195
rect 35345 6125 35415 6155
rect 36545 6195 36615 6210
rect 36545 6155 36560 6195
rect 36600 6155 36615 6195
rect 36545 6125 36615 6155
rect 37025 6195 37095 6210
rect 37025 6155 37040 6195
rect 37080 6155 37095 6195
rect 37025 6125 37095 6155
rect 38225 6195 38295 6210
rect 38225 6155 38240 6195
rect 38280 6155 38295 6195
rect 38225 6125 38295 6155
rect 40300 6195 40370 6210
rect 40300 6155 40315 6195
rect 40355 6155 40370 6195
rect 40300 6125 40370 6155
rect 41500 6195 41570 6210
rect 41500 6155 41515 6195
rect 41555 6155 41570 6195
rect 41500 6125 41570 6155
rect 41980 6195 42050 6210
rect 41980 6155 41995 6195
rect 42035 6155 42050 6195
rect 41980 6125 42050 6155
rect 43180 6195 43250 6210
rect 43180 6155 43195 6195
rect 43235 6155 43250 6195
rect 43180 6125 43250 6155
rect 45255 6195 45325 6210
rect 45255 6155 45270 6195
rect 45310 6155 45325 6195
rect 45255 6125 45325 6155
rect 46455 6195 46525 6210
rect 46455 6155 46470 6195
rect 46510 6155 46525 6195
rect 46455 6125 46525 6155
rect 46935 6195 47005 6210
rect 46935 6155 46950 6195
rect 46990 6155 47005 6195
rect 46935 6125 47005 6155
rect 48135 6195 48205 6210
rect 48135 6155 48150 6195
rect 48190 6155 48205 6195
rect 48135 6125 48205 6155
rect 50210 6195 50280 6210
rect 50210 6155 50225 6195
rect 50265 6155 50280 6195
rect 50210 6125 50280 6155
rect 51410 6195 51480 6210
rect 51410 6155 51425 6195
rect 51465 6155 51480 6195
rect 51410 6125 51480 6155
rect 51890 6195 51960 6210
rect 51890 6155 51905 6195
rect 51945 6155 51960 6195
rect 51890 6125 51960 6155
rect 53090 6195 53160 6210
rect 53090 6155 53105 6195
rect 53145 6155 53160 6195
rect 53090 6125 53160 6155
rect 55165 6195 55235 6210
rect 55165 6155 55180 6195
rect 55220 6155 55235 6195
rect 55165 6125 55235 6155
rect 56365 6195 56435 6210
rect 56365 6155 56380 6195
rect 56420 6155 56435 6195
rect 56365 6125 56435 6155
rect 56845 6195 56915 6210
rect 56845 6155 56860 6195
rect 56900 6155 56915 6195
rect 56845 6125 56915 6155
rect 58045 6195 58115 6210
rect 58045 6155 58060 6195
rect 58100 6155 58115 6195
rect 58045 6125 58115 6155
rect 60120 6195 60190 6210
rect 60120 6155 60135 6195
rect 60175 6155 60190 6195
rect 60120 6125 60190 6155
rect 61320 6195 61390 6210
rect 61320 6155 61335 6195
rect 61375 6155 61390 6195
rect 61320 6125 61390 6155
rect 61800 6195 61870 6210
rect 61800 6155 61815 6195
rect 61855 6155 61870 6195
rect 61800 6125 61870 6155
rect 63000 6195 63070 6210
rect 63000 6155 63015 6195
rect 63055 6155 63070 6195
rect 63000 6125 63070 6155
rect 65075 6195 65145 6210
rect 65075 6155 65090 6195
rect 65130 6155 65145 6195
rect 65075 6125 65145 6155
rect 66275 6195 66345 6210
rect 66275 6155 66290 6195
rect 66330 6155 66345 6195
rect 66275 6125 66345 6155
rect 66755 6195 66825 6210
rect 66755 6155 66770 6195
rect 66810 6155 66825 6195
rect 66755 6125 66825 6155
rect 67955 6195 68025 6210
rect 67955 6155 67970 6195
rect 68010 6155 68025 6195
rect 67955 6125 68025 6155
rect 70030 6195 70100 6210
rect 70030 6155 70045 6195
rect 70085 6155 70100 6195
rect 70030 6125 70100 6155
rect 71230 6195 71300 6210
rect 71230 6155 71245 6195
rect 71285 6155 71300 6195
rect 71230 6125 71300 6155
rect 71710 6195 71780 6210
rect 71710 6155 71725 6195
rect 71765 6155 71780 6195
rect 71710 6125 71780 6155
rect 72910 6195 72980 6210
rect 72910 6155 72925 6195
rect 72965 6155 72980 6195
rect 72910 6125 72980 6155
rect 74985 6195 75055 6210
rect 74985 6155 75000 6195
rect 75040 6155 75055 6195
rect 74985 6125 75055 6155
rect 76185 6195 76255 6210
rect 76185 6155 76200 6195
rect 76240 6155 76255 6195
rect 76185 6125 76255 6155
rect 76665 6195 76735 6210
rect 76665 6155 76680 6195
rect 76720 6155 76735 6195
rect 76665 6125 76735 6155
rect 77865 6195 77935 6210
rect 77865 6155 77880 6195
rect 77920 6155 77935 6195
rect 77865 6125 77935 6155
rect 660 5885 77935 5900
rect 660 5850 675 5885
rect 715 5850 1875 5885
rect 1915 5850 2355 5885
rect 2395 5850 3555 5885
rect 3595 5850 5630 5885
rect 5670 5850 6830 5885
rect 6870 5850 7310 5885
rect 7350 5850 8510 5885
rect 8550 5850 10585 5885
rect 10625 5850 11785 5885
rect 11825 5850 12265 5885
rect 12305 5850 13465 5885
rect 13505 5850 15540 5885
rect 15580 5850 16740 5885
rect 16780 5850 17220 5885
rect 17260 5850 18420 5885
rect 18460 5850 20495 5885
rect 20535 5850 21695 5885
rect 21735 5850 22175 5885
rect 22215 5850 23375 5885
rect 23415 5850 25450 5885
rect 25490 5850 26650 5885
rect 26690 5850 27130 5885
rect 27170 5850 28330 5885
rect 28370 5850 30405 5885
rect 30445 5850 31605 5885
rect 31645 5850 32085 5885
rect 32125 5850 33285 5885
rect 33325 5850 35360 5885
rect 35400 5850 36560 5885
rect 36600 5850 37040 5885
rect 37080 5850 38240 5885
rect 38280 5850 40315 5885
rect 40355 5850 41515 5885
rect 41555 5850 41995 5885
rect 42035 5850 43195 5885
rect 43235 5850 45270 5885
rect 45310 5850 46470 5885
rect 46510 5850 46950 5885
rect 46990 5850 48150 5885
rect 48190 5850 50225 5885
rect 50265 5850 51425 5885
rect 51465 5850 51905 5885
rect 51945 5850 53105 5885
rect 53145 5850 55180 5885
rect 55220 5850 56380 5885
rect 56420 5850 56860 5885
rect 56900 5850 58060 5885
rect 58100 5850 60135 5885
rect 60175 5850 61335 5885
rect 61375 5850 61815 5885
rect 61855 5850 63015 5885
rect 63055 5850 65090 5885
rect 65130 5850 66290 5885
rect 66330 5850 66770 5885
rect 66810 5850 67970 5885
rect 68010 5850 70045 5885
rect 70085 5850 71245 5885
rect 71285 5850 71725 5885
rect 71765 5850 72925 5885
rect 72965 5850 75000 5885
rect 75040 5850 76200 5885
rect 76240 5850 76680 5885
rect 76720 5850 77880 5885
rect 77920 5850 77935 5885
rect 660 5835 77935 5850
rect 5615 5565 5685 5595
rect 5615 5525 5630 5565
rect 5670 5525 5685 5565
rect 5615 5510 5685 5525
rect 6815 5565 6885 5595
rect 6815 5525 6830 5565
rect 6870 5525 6885 5565
rect 6815 5510 6885 5525
rect 7295 5565 7365 5595
rect 7295 5525 7310 5565
rect 7350 5525 7365 5565
rect 7295 5510 7365 5525
rect 8495 5565 8565 5595
rect 8495 5525 8510 5565
rect 8550 5525 8565 5565
rect 8495 5510 8565 5525
rect 10570 5565 10640 5595
rect 10570 5525 10585 5565
rect 10625 5525 10640 5565
rect 10570 5510 10640 5525
rect 11770 5565 11840 5595
rect 11770 5525 11785 5565
rect 11825 5525 11840 5565
rect 11770 5510 11840 5525
rect 12250 5565 12320 5595
rect 12250 5525 12265 5565
rect 12305 5525 12320 5565
rect 12250 5510 12320 5525
rect 13450 5565 13520 5595
rect 13450 5525 13465 5565
rect 13505 5525 13520 5565
rect 13450 5510 13520 5525
rect 15525 5565 15595 5595
rect 15525 5525 15540 5565
rect 15580 5525 15595 5565
rect 15525 5510 15595 5525
rect 16725 5565 16795 5595
rect 16725 5525 16740 5565
rect 16780 5525 16795 5565
rect 16725 5510 16795 5525
rect 17205 5565 17275 5595
rect 17205 5525 17220 5565
rect 17260 5525 17275 5565
rect 17205 5510 17275 5525
rect 18405 5565 18475 5595
rect 18405 5525 18420 5565
rect 18460 5525 18475 5565
rect 18405 5510 18475 5525
rect 20480 5565 20550 5595
rect 20480 5525 20495 5565
rect 20535 5525 20550 5565
rect 20480 5510 20550 5525
rect 21680 5565 21750 5595
rect 21680 5525 21695 5565
rect 21735 5525 21750 5565
rect 21680 5510 21750 5525
rect 22160 5565 22230 5595
rect 22160 5525 22175 5565
rect 22215 5525 22230 5565
rect 22160 5510 22230 5525
rect 23360 5565 23430 5595
rect 23360 5525 23375 5565
rect 23415 5525 23430 5565
rect 23360 5510 23430 5525
rect 25435 5565 25505 5595
rect 25435 5525 25450 5565
rect 25490 5525 25505 5565
rect 25435 5510 25505 5525
rect 26635 5565 26705 5595
rect 26635 5525 26650 5565
rect 26690 5525 26705 5565
rect 26635 5510 26705 5525
rect 27115 5565 27185 5595
rect 27115 5525 27130 5565
rect 27170 5525 27185 5565
rect 27115 5510 27185 5525
rect 28315 5565 28385 5595
rect 28315 5525 28330 5565
rect 28370 5525 28385 5565
rect 28315 5510 28385 5525
rect 30390 5565 30460 5595
rect 30390 5525 30405 5565
rect 30445 5525 30460 5565
rect 30390 5510 30460 5525
rect 31590 5565 31660 5595
rect 31590 5525 31605 5565
rect 31645 5525 31660 5565
rect 31590 5510 31660 5525
rect 32070 5565 32140 5595
rect 32070 5525 32085 5565
rect 32125 5525 32140 5565
rect 32070 5510 32140 5525
rect 33270 5565 33340 5595
rect 33270 5525 33285 5565
rect 33325 5525 33340 5565
rect 33270 5510 33340 5525
rect 35345 5565 35415 5595
rect 35345 5525 35360 5565
rect 35400 5525 35415 5565
rect 35345 5510 35415 5525
rect 36545 5565 36615 5595
rect 36545 5525 36560 5565
rect 36600 5525 36615 5565
rect 36545 5510 36615 5525
rect 37025 5565 37095 5595
rect 37025 5525 37040 5565
rect 37080 5525 37095 5565
rect 37025 5510 37095 5525
rect 38225 5565 38295 5595
rect 38225 5525 38240 5565
rect 38280 5525 38295 5565
rect 38225 5510 38295 5525
rect 40300 5565 40370 5595
rect 40300 5525 40315 5565
rect 40355 5525 40370 5565
rect 40300 5510 40370 5525
rect 41500 5565 41570 5595
rect 41500 5525 41515 5565
rect 41555 5525 41570 5565
rect 41500 5510 41570 5525
rect 41980 5565 42050 5595
rect 41980 5525 41995 5565
rect 42035 5525 42050 5565
rect 41980 5510 42050 5525
rect 43180 5565 43250 5595
rect 43180 5525 43195 5565
rect 43235 5525 43250 5565
rect 43180 5510 43250 5525
rect 45255 5565 45325 5595
rect 45255 5525 45270 5565
rect 45310 5525 45325 5565
rect 45255 5510 45325 5525
rect 46455 5565 46525 5595
rect 46455 5525 46470 5565
rect 46510 5525 46525 5565
rect 46455 5510 46525 5525
rect 46935 5565 47005 5595
rect 46935 5525 46950 5565
rect 46990 5525 47005 5565
rect 46935 5510 47005 5525
rect 48135 5565 48205 5595
rect 48135 5525 48150 5565
rect 48190 5525 48205 5565
rect 48135 5510 48205 5525
rect 50210 5565 50280 5595
rect 50210 5525 50225 5565
rect 50265 5525 50280 5565
rect 50210 5510 50280 5525
rect 51410 5565 51480 5595
rect 51410 5525 51425 5565
rect 51465 5525 51480 5565
rect 51410 5510 51480 5525
rect 51890 5565 51960 5595
rect 51890 5525 51905 5565
rect 51945 5525 51960 5565
rect 51890 5510 51960 5525
rect 53090 5565 53160 5595
rect 53090 5525 53105 5565
rect 53145 5525 53160 5565
rect 53090 5510 53160 5525
rect 55165 5565 55235 5595
rect 55165 5525 55180 5565
rect 55220 5525 55235 5565
rect 55165 5510 55235 5525
rect 56365 5565 56435 5595
rect 56365 5525 56380 5565
rect 56420 5525 56435 5565
rect 56365 5510 56435 5525
rect 56845 5565 56915 5595
rect 56845 5525 56860 5565
rect 56900 5525 56915 5565
rect 56845 5510 56915 5525
rect 58045 5565 58115 5595
rect 58045 5525 58060 5565
rect 58100 5525 58115 5565
rect 58045 5510 58115 5525
rect 60120 5565 60190 5595
rect 60120 5525 60135 5565
rect 60175 5525 60190 5565
rect 60120 5510 60190 5525
rect 61320 5565 61390 5595
rect 61320 5525 61335 5565
rect 61375 5525 61390 5565
rect 61320 5510 61390 5525
rect 61800 5565 61870 5595
rect 61800 5525 61815 5565
rect 61855 5525 61870 5565
rect 61800 5510 61870 5525
rect 63000 5565 63070 5595
rect 63000 5525 63015 5565
rect 63055 5525 63070 5565
rect 63000 5510 63070 5525
rect 65075 5565 65145 5595
rect 65075 5525 65090 5565
rect 65130 5525 65145 5565
rect 65075 5510 65145 5525
rect 66275 5565 66345 5595
rect 66275 5525 66290 5565
rect 66330 5525 66345 5565
rect 66275 5510 66345 5525
rect 66755 5565 66825 5595
rect 66755 5525 66770 5565
rect 66810 5525 66825 5565
rect 66755 5510 66825 5525
rect 67955 5565 68025 5595
rect 67955 5525 67970 5565
rect 68010 5525 68025 5565
rect 67955 5510 68025 5525
rect 70030 5565 70100 5595
rect 70030 5525 70045 5565
rect 70085 5525 70100 5565
rect 70030 5510 70100 5525
rect 71230 5565 71300 5595
rect 71230 5525 71245 5565
rect 71285 5525 71300 5565
rect 71230 5510 71300 5525
rect 71710 5565 71780 5595
rect 71710 5525 71725 5565
rect 71765 5525 71780 5565
rect 71710 5510 71780 5525
rect 72910 5565 72980 5595
rect 72910 5525 72925 5565
rect 72965 5525 72980 5565
rect 72910 5510 72980 5525
rect 74985 5565 75055 5595
rect 74985 5525 75000 5565
rect 75040 5525 75055 5565
rect 74985 5510 75055 5525
rect 76185 5565 76255 5595
rect 76185 5525 76200 5565
rect 76240 5525 76255 5565
rect 76185 5510 76255 5525
rect 76665 5565 76735 5595
rect 76665 5525 76680 5565
rect 76720 5525 76735 5565
rect 76665 5510 76735 5525
rect 77865 5565 77935 5595
rect 77865 5525 77880 5565
rect 77920 5525 77935 5565
rect 77865 5510 77935 5525
rect -345 5480 -280 5495
rect -345 5445 -330 5480
rect -295 5460 -280 5480
rect -295 5445 0 5460
rect -345 5430 0 5445
rect 4295 5430 4955 5460
rect 9250 5430 9910 5460
rect 14205 5430 14865 5460
rect 19160 5430 19820 5460
rect 24115 5430 24775 5460
rect 29070 5430 29730 5460
rect 34025 5430 34685 5460
rect 38980 5430 39640 5460
rect 43935 5430 44595 5460
rect 48890 5430 49550 5460
rect 53845 5430 54505 5460
rect 58800 5430 59460 5460
rect 63755 5430 64415 5460
rect 68710 5430 69370 5460
rect 73665 5430 74325 5460
rect 8690 5325 8775 5340
rect 8690 5285 8705 5325
rect 8745 5285 8775 5325
rect 8690 5270 8775 5285
rect 10355 5325 10440 5340
rect 10355 5285 10385 5325
rect 10425 5285 10440 5325
rect 10355 5270 10440 5285
rect 13645 5325 13730 5340
rect 13645 5285 13660 5325
rect 13700 5285 13730 5325
rect 13645 5270 13730 5285
rect 15310 5325 15395 5340
rect 15310 5285 15340 5325
rect 15380 5285 15395 5325
rect 15310 5270 15395 5285
rect 18600 5325 18685 5340
rect 18600 5285 18615 5325
rect 18655 5285 18685 5325
rect 18600 5270 18685 5285
rect 20265 5325 20350 5340
rect 20265 5285 20295 5325
rect 20335 5285 20350 5325
rect 20265 5270 20350 5285
rect 23555 5325 23640 5340
rect 23555 5285 23570 5325
rect 23610 5285 23640 5325
rect 23555 5270 23640 5285
rect 25220 5325 25305 5340
rect 25220 5285 25250 5325
rect 25290 5285 25305 5325
rect 25220 5270 25305 5285
rect 28510 5325 28595 5340
rect 28510 5285 28525 5325
rect 28565 5285 28595 5325
rect 28510 5270 28595 5285
rect 30175 5325 30260 5340
rect 30175 5285 30205 5325
rect 30245 5285 30260 5325
rect 30175 5270 30260 5285
rect 33465 5325 33550 5340
rect 33465 5285 33480 5325
rect 33520 5285 33550 5325
rect 33465 5270 33550 5285
rect 35130 5325 35215 5340
rect 35130 5285 35160 5325
rect 35200 5285 35215 5325
rect 35130 5270 35215 5285
rect 38420 5325 38505 5340
rect 38420 5285 38435 5325
rect 38475 5285 38505 5325
rect 38420 5270 38505 5285
rect 40085 5325 40170 5340
rect 40085 5285 40115 5325
rect 40155 5285 40170 5325
rect 40085 5270 40170 5285
rect 43375 5325 43460 5340
rect 43375 5285 43390 5325
rect 43430 5285 43460 5325
rect 43375 5270 43460 5285
rect 45040 5325 45125 5340
rect 45040 5285 45070 5325
rect 45110 5285 45125 5325
rect 45040 5270 45125 5285
rect 48330 5325 48415 5340
rect 48330 5285 48345 5325
rect 48385 5285 48415 5325
rect 48330 5270 48415 5285
rect 49995 5325 50080 5340
rect 49995 5285 50025 5325
rect 50065 5285 50080 5325
rect 49995 5270 50080 5285
rect 53285 5325 53370 5340
rect 53285 5285 53300 5325
rect 53340 5285 53370 5325
rect 53285 5270 53370 5285
rect 54950 5325 55035 5340
rect 54950 5285 54980 5325
rect 55020 5285 55035 5325
rect 54950 5270 55035 5285
rect 58240 5325 58325 5340
rect 58240 5285 58255 5325
rect 58295 5285 58325 5325
rect 58240 5270 58325 5285
rect 59905 5325 59990 5340
rect 59905 5285 59935 5325
rect 59975 5285 59990 5325
rect 59905 5270 59990 5285
rect 63195 5325 63280 5340
rect 63195 5285 63210 5325
rect 63250 5285 63280 5325
rect 63195 5270 63280 5285
rect 64860 5325 64945 5340
rect 64860 5285 64890 5325
rect 64930 5285 64945 5325
rect 64860 5270 64945 5285
rect 68150 5325 68235 5340
rect 68150 5285 68165 5325
rect 68205 5285 68235 5325
rect 68150 5270 68235 5285
rect 69815 5325 69900 5340
rect 69815 5285 69845 5325
rect 69885 5285 69900 5325
rect 69815 5270 69900 5285
rect 73105 5325 73190 5340
rect 73105 5285 73120 5325
rect 73160 5285 73190 5325
rect 73105 5270 73190 5285
rect 74770 5325 74855 5340
rect 74770 5285 74800 5325
rect 74840 5285 74855 5325
rect 74770 5270 74855 5285
rect 8690 3405 8775 3420
rect 8690 3365 8705 3405
rect 8745 3365 8775 3405
rect 8690 3350 8775 3365
rect 10355 3405 10440 3420
rect 10355 3365 10385 3405
rect 10425 3365 10440 3405
rect 10355 3350 10440 3365
rect 13645 3405 13730 3420
rect 13645 3365 13660 3405
rect 13700 3365 13730 3405
rect 13645 3350 13730 3365
rect 15310 3405 15395 3420
rect 15310 3365 15340 3405
rect 15380 3365 15395 3405
rect 15310 3350 15395 3365
rect 18600 3405 18685 3420
rect 18600 3365 18615 3405
rect 18655 3365 18685 3405
rect 18600 3350 18685 3365
rect 20265 3405 20350 3420
rect 20265 3365 20295 3405
rect 20335 3365 20350 3405
rect 20265 3350 20350 3365
rect 23555 3405 23640 3420
rect 23555 3365 23570 3405
rect 23610 3365 23640 3405
rect 23555 3350 23640 3365
rect 25220 3405 25305 3420
rect 25220 3365 25250 3405
rect 25290 3365 25305 3405
rect 25220 3350 25305 3365
rect 28510 3405 28595 3420
rect 28510 3365 28525 3405
rect 28565 3365 28595 3405
rect 28510 3350 28595 3365
rect 30175 3405 30260 3420
rect 30175 3365 30205 3405
rect 30245 3365 30260 3405
rect 30175 3350 30260 3365
rect 33465 3405 33550 3420
rect 33465 3365 33480 3405
rect 33520 3365 33550 3405
rect 33465 3350 33550 3365
rect 35130 3405 35215 3420
rect 35130 3365 35160 3405
rect 35200 3365 35215 3405
rect 35130 3350 35215 3365
rect 38420 3405 38505 3420
rect 38420 3365 38435 3405
rect 38475 3365 38505 3405
rect 38420 3350 38505 3365
rect 40085 3405 40170 3420
rect 40085 3365 40115 3405
rect 40155 3365 40170 3405
rect 40085 3350 40170 3365
rect 43375 3405 43460 3420
rect 43375 3365 43390 3405
rect 43430 3365 43460 3405
rect 43375 3350 43460 3365
rect 45040 3405 45125 3420
rect 45040 3365 45070 3405
rect 45110 3365 45125 3405
rect 45040 3350 45125 3365
rect 48330 3405 48415 3420
rect 48330 3365 48345 3405
rect 48385 3365 48415 3405
rect 48330 3350 48415 3365
rect 49995 3405 50080 3420
rect 49995 3365 50025 3405
rect 50065 3365 50080 3405
rect 49995 3350 50080 3365
rect 53285 3405 53370 3420
rect 53285 3365 53300 3405
rect 53340 3365 53370 3405
rect 53285 3350 53370 3365
rect 54950 3405 55035 3420
rect 54950 3365 54980 3405
rect 55020 3365 55035 3405
rect 54950 3350 55035 3365
rect 58240 3405 58325 3420
rect 58240 3365 58255 3405
rect 58295 3365 58325 3405
rect 58240 3350 58325 3365
rect 59905 3405 59990 3420
rect 59905 3365 59935 3405
rect 59975 3365 59990 3405
rect 59905 3350 59990 3365
rect 63195 3405 63280 3420
rect 63195 3365 63210 3405
rect 63250 3365 63280 3405
rect 63195 3350 63280 3365
rect 64860 3405 64945 3420
rect 64860 3365 64890 3405
rect 64930 3365 64945 3405
rect 64860 3350 64945 3365
rect 68150 3405 68235 3420
rect 68150 3365 68165 3405
rect 68205 3365 68235 3405
rect 68150 3350 68235 3365
rect 69815 3405 69900 3420
rect 69815 3365 69845 3405
rect 69885 3365 69900 3405
rect 69815 3350 69900 3365
rect 73105 3405 73190 3420
rect 73105 3365 73120 3405
rect 73160 3365 73190 3405
rect 73105 3350 73190 3365
rect 74770 3405 74855 3420
rect 74770 3365 74800 3405
rect 74840 3365 74855 3405
rect 74770 3350 74855 3365
rect 15 3260 80 3275
rect 15 3225 30 3260
rect 65 3225 80 3260
rect 15 3210 80 3225
rect 4365 3210 4970 3240
rect 9320 3210 9925 3240
rect 14275 3210 14880 3240
rect 19230 3210 19835 3240
rect 24185 3210 24790 3240
rect 29140 3210 29745 3240
rect 34095 3210 34700 3240
rect 39050 3210 39655 3240
rect 44005 3210 44610 3240
rect 48960 3210 49565 3240
rect 53915 3210 54520 3240
rect 58870 3210 59475 3240
rect 63825 3210 64430 3240
rect 68780 3210 69385 3240
rect 73735 3210 74340 3240
rect 660 3120 730 3135
rect 660 3080 675 3120
rect 715 3080 730 3120
rect 660 3050 730 3080
rect 5615 3120 5685 3135
rect 5615 3080 5630 3120
rect 5670 3080 5685 3120
rect 5615 3050 5685 3080
rect 6815 3120 6885 3135
rect 6815 3080 6830 3120
rect 6870 3080 6885 3120
rect 6815 3050 6885 3080
rect 7295 3120 7365 3135
rect 7295 3080 7310 3120
rect 7350 3080 7365 3120
rect 7295 3050 7365 3080
rect 8495 3120 8565 3135
rect 8495 3080 8510 3120
rect 8550 3080 8565 3120
rect 8495 3050 8565 3080
rect 10570 3120 10640 3135
rect 10570 3080 10585 3120
rect 10625 3080 10640 3120
rect 10570 3050 10640 3080
rect 11770 3120 11840 3135
rect 11770 3080 11785 3120
rect 11825 3080 11840 3120
rect 11770 3050 11840 3080
rect 12250 3120 12320 3135
rect 12250 3080 12265 3120
rect 12305 3080 12320 3120
rect 12250 3050 12320 3080
rect 13450 3120 13520 3135
rect 13450 3080 13465 3120
rect 13505 3080 13520 3120
rect 13450 3050 13520 3080
rect 15525 3120 15595 3135
rect 15525 3080 15540 3120
rect 15580 3080 15595 3120
rect 15525 3050 15595 3080
rect 16725 3120 16795 3135
rect 16725 3080 16740 3120
rect 16780 3080 16795 3120
rect 16725 3050 16795 3080
rect 17205 3120 17275 3135
rect 17205 3080 17220 3120
rect 17260 3080 17275 3120
rect 17205 3050 17275 3080
rect 18405 3120 18475 3135
rect 18405 3080 18420 3120
rect 18460 3080 18475 3120
rect 18405 3050 18475 3080
rect 20480 3120 20550 3135
rect 20480 3080 20495 3120
rect 20535 3080 20550 3120
rect 20480 3050 20550 3080
rect 21680 3120 21750 3135
rect 21680 3080 21695 3120
rect 21735 3080 21750 3120
rect 21680 3050 21750 3080
rect 22160 3120 22230 3135
rect 22160 3080 22175 3120
rect 22215 3080 22230 3120
rect 22160 3050 22230 3080
rect 23360 3120 23430 3135
rect 23360 3080 23375 3120
rect 23415 3080 23430 3120
rect 23360 3050 23430 3080
rect 25435 3120 25505 3135
rect 25435 3080 25450 3120
rect 25490 3080 25505 3120
rect 25435 3050 25505 3080
rect 26635 3120 26705 3135
rect 26635 3080 26650 3120
rect 26690 3080 26705 3120
rect 26635 3050 26705 3080
rect 27115 3120 27185 3135
rect 27115 3080 27130 3120
rect 27170 3080 27185 3120
rect 27115 3050 27185 3080
rect 28315 3120 28385 3135
rect 28315 3080 28330 3120
rect 28370 3080 28385 3120
rect 28315 3050 28385 3080
rect 30390 3120 30460 3135
rect 30390 3080 30405 3120
rect 30445 3080 30460 3120
rect 30390 3050 30460 3080
rect 31590 3120 31660 3135
rect 31590 3080 31605 3120
rect 31645 3080 31660 3120
rect 31590 3050 31660 3080
rect 32070 3120 32140 3135
rect 32070 3080 32085 3120
rect 32125 3080 32140 3120
rect 32070 3050 32140 3080
rect 33270 3120 33340 3135
rect 33270 3080 33285 3120
rect 33325 3080 33340 3120
rect 33270 3050 33340 3080
rect 35345 3120 35415 3135
rect 35345 3080 35360 3120
rect 35400 3080 35415 3120
rect 35345 3050 35415 3080
rect 36545 3120 36615 3135
rect 36545 3080 36560 3120
rect 36600 3080 36615 3120
rect 36545 3050 36615 3080
rect 37025 3120 37095 3135
rect 37025 3080 37040 3120
rect 37080 3080 37095 3120
rect 37025 3050 37095 3080
rect 38225 3120 38295 3135
rect 38225 3080 38240 3120
rect 38280 3080 38295 3120
rect 38225 3050 38295 3080
rect 40300 3120 40370 3135
rect 40300 3080 40315 3120
rect 40355 3080 40370 3120
rect 40300 3050 40370 3080
rect 41500 3120 41570 3135
rect 41500 3080 41515 3120
rect 41555 3080 41570 3120
rect 41500 3050 41570 3080
rect 41980 3120 42050 3135
rect 41980 3080 41995 3120
rect 42035 3080 42050 3120
rect 41980 3050 42050 3080
rect 43180 3120 43250 3135
rect 43180 3080 43195 3120
rect 43235 3080 43250 3120
rect 43180 3050 43250 3080
rect 45255 3120 45325 3135
rect 45255 3080 45270 3120
rect 45310 3080 45325 3120
rect 45255 3050 45325 3080
rect 46455 3120 46525 3135
rect 46455 3080 46470 3120
rect 46510 3080 46525 3120
rect 46455 3050 46525 3080
rect 46935 3120 47005 3135
rect 46935 3080 46950 3120
rect 46990 3080 47005 3120
rect 46935 3050 47005 3080
rect 48135 3120 48205 3135
rect 48135 3080 48150 3120
rect 48190 3080 48205 3120
rect 48135 3050 48205 3080
rect 50210 3120 50280 3135
rect 50210 3080 50225 3120
rect 50265 3080 50280 3120
rect 50210 3050 50280 3080
rect 51410 3120 51480 3135
rect 51410 3080 51425 3120
rect 51465 3080 51480 3120
rect 51410 3050 51480 3080
rect 51890 3120 51960 3135
rect 51890 3080 51905 3120
rect 51945 3080 51960 3120
rect 51890 3050 51960 3080
rect 53090 3120 53160 3135
rect 53090 3080 53105 3120
rect 53145 3080 53160 3120
rect 53090 3050 53160 3080
rect 55165 3120 55235 3135
rect 55165 3080 55180 3120
rect 55220 3080 55235 3120
rect 55165 3050 55235 3080
rect 56365 3120 56435 3135
rect 56365 3080 56380 3120
rect 56420 3080 56435 3120
rect 56365 3050 56435 3080
rect 56845 3120 56915 3135
rect 56845 3080 56860 3120
rect 56900 3080 56915 3120
rect 56845 3050 56915 3080
rect 58045 3120 58115 3135
rect 58045 3080 58060 3120
rect 58100 3080 58115 3120
rect 58045 3050 58115 3080
rect 60120 3120 60190 3135
rect 60120 3080 60135 3120
rect 60175 3080 60190 3120
rect 60120 3050 60190 3080
rect 61320 3120 61390 3135
rect 61320 3080 61335 3120
rect 61375 3080 61390 3120
rect 61320 3050 61390 3080
rect 61800 3120 61870 3135
rect 61800 3080 61815 3120
rect 61855 3080 61870 3120
rect 61800 3050 61870 3080
rect 63000 3120 63070 3135
rect 63000 3080 63015 3120
rect 63055 3080 63070 3120
rect 63000 3050 63070 3080
rect 65075 3120 65145 3135
rect 65075 3080 65090 3120
rect 65130 3080 65145 3120
rect 65075 3050 65145 3080
rect 66275 3120 66345 3135
rect 66275 3080 66290 3120
rect 66330 3080 66345 3120
rect 66275 3050 66345 3080
rect 66755 3120 66825 3135
rect 66755 3080 66770 3120
rect 66810 3080 66825 3120
rect 66755 3050 66825 3080
rect 67955 3120 68025 3135
rect 67955 3080 67970 3120
rect 68010 3080 68025 3120
rect 67955 3050 68025 3080
rect 70030 3120 70100 3135
rect 70030 3080 70045 3120
rect 70085 3080 70100 3120
rect 70030 3050 70100 3080
rect 71230 3120 71300 3135
rect 71230 3080 71245 3120
rect 71285 3080 71300 3120
rect 71230 3050 71300 3080
rect 71710 3120 71780 3135
rect 71710 3080 71725 3120
rect 71765 3080 71780 3120
rect 71710 3050 71780 3080
rect 72910 3120 72980 3135
rect 72910 3080 72925 3120
rect 72965 3080 72980 3120
rect 72910 3050 72980 3080
rect 74985 3120 75055 3135
rect 74985 3080 75000 3120
rect 75040 3080 75055 3120
rect 74985 3050 75055 3080
rect 76185 3120 76255 3135
rect 76185 3080 76200 3120
rect 76240 3080 76255 3120
rect 76185 3050 76255 3080
rect 76665 3120 76735 3135
rect 76665 3080 76680 3120
rect 76720 3080 76735 3120
rect 76665 3050 76735 3080
rect 77865 3120 77935 3135
rect 77865 3080 77880 3120
rect 77920 3080 77935 3120
rect 77865 3050 77935 3080
rect 660 2835 77935 2850
rect 660 2800 675 2835
rect 715 2800 1875 2835
rect 1915 2800 2355 2835
rect 2395 2800 3555 2835
rect 3595 2800 5630 2835
rect 5670 2800 6830 2835
rect 6870 2800 7310 2835
rect 7350 2800 8510 2835
rect 8550 2800 10585 2835
rect 10625 2800 11785 2835
rect 11825 2800 12265 2835
rect 12305 2800 13465 2835
rect 13505 2800 15540 2835
rect 15580 2800 16740 2835
rect 16780 2800 17220 2835
rect 17260 2800 18420 2835
rect 18460 2800 20495 2835
rect 20535 2800 21695 2835
rect 21735 2800 22175 2835
rect 22215 2800 23375 2835
rect 23415 2800 25450 2835
rect 25490 2800 26650 2835
rect 26690 2800 27130 2835
rect 27170 2800 28330 2835
rect 28370 2800 30405 2835
rect 30445 2800 31605 2835
rect 31645 2800 32085 2835
rect 32125 2800 33285 2835
rect 33325 2800 35360 2835
rect 35400 2800 36560 2835
rect 36600 2800 37040 2835
rect 37080 2800 38240 2835
rect 38280 2800 40315 2835
rect 40355 2800 41515 2835
rect 41555 2800 41995 2835
rect 42035 2800 43195 2835
rect 43235 2800 45270 2835
rect 45310 2800 46470 2835
rect 46510 2800 46950 2835
rect 46990 2800 48150 2835
rect 48190 2800 50225 2835
rect 50265 2800 51425 2835
rect 51465 2800 51905 2835
rect 51945 2800 53105 2835
rect 53145 2800 55180 2835
rect 55220 2800 56380 2835
rect 56420 2800 56860 2835
rect 56900 2800 58060 2835
rect 58100 2800 60135 2835
rect 60175 2800 61335 2835
rect 61375 2800 61815 2835
rect 61855 2800 63015 2835
rect 63055 2800 65090 2835
rect 65130 2800 66290 2835
rect 66330 2800 66770 2835
rect 66810 2800 67970 2835
rect 68010 2800 70045 2835
rect 70085 2800 71245 2835
rect 71285 2800 71725 2835
rect 71765 2800 72925 2835
rect 72965 2800 75000 2835
rect 75040 2800 76200 2835
rect 76240 2800 76680 2835
rect 76720 2800 77880 2835
rect 77920 2800 77935 2835
rect 660 2785 77935 2800
rect 660 2490 730 2520
rect 660 2450 675 2490
rect 715 2450 730 2490
rect 660 2435 730 2450
rect 5615 2490 5685 2520
rect 5615 2450 5630 2490
rect 5670 2450 5685 2490
rect 5615 2435 5685 2450
rect 6815 2490 6885 2520
rect 6815 2450 6830 2490
rect 6870 2450 6885 2490
rect 6815 2435 6885 2450
rect 7295 2490 7365 2520
rect 7295 2450 7310 2490
rect 7350 2450 7365 2490
rect 7295 2435 7365 2450
rect 8495 2490 8565 2520
rect 8495 2450 8510 2490
rect 8550 2450 8565 2490
rect 8495 2435 8565 2450
rect 10570 2490 10640 2520
rect 10570 2450 10585 2490
rect 10625 2450 10640 2490
rect 10570 2435 10640 2450
rect 11770 2490 11840 2520
rect 11770 2450 11785 2490
rect 11825 2450 11840 2490
rect 11770 2435 11840 2450
rect 12250 2490 12320 2520
rect 12250 2450 12265 2490
rect 12305 2450 12320 2490
rect 12250 2435 12320 2450
rect 13450 2490 13520 2520
rect 13450 2450 13465 2490
rect 13505 2450 13520 2490
rect 13450 2435 13520 2450
rect 15525 2490 15595 2520
rect 15525 2450 15540 2490
rect 15580 2450 15595 2490
rect 15525 2435 15595 2450
rect 16725 2490 16795 2520
rect 16725 2450 16740 2490
rect 16780 2450 16795 2490
rect 16725 2435 16795 2450
rect 17205 2490 17275 2520
rect 17205 2450 17220 2490
rect 17260 2450 17275 2490
rect 17205 2435 17275 2450
rect 18405 2490 18475 2520
rect 18405 2450 18420 2490
rect 18460 2450 18475 2490
rect 18405 2435 18475 2450
rect 20480 2490 20550 2520
rect 20480 2450 20495 2490
rect 20535 2450 20550 2490
rect 20480 2435 20550 2450
rect 21680 2490 21750 2520
rect 21680 2450 21695 2490
rect 21735 2450 21750 2490
rect 21680 2435 21750 2450
rect 22160 2490 22230 2520
rect 22160 2450 22175 2490
rect 22215 2450 22230 2490
rect 22160 2435 22230 2450
rect 23360 2490 23430 2520
rect 23360 2450 23375 2490
rect 23415 2450 23430 2490
rect 23360 2435 23430 2450
rect 25435 2490 25505 2520
rect 25435 2450 25450 2490
rect 25490 2450 25505 2490
rect 25435 2435 25505 2450
rect 26635 2490 26705 2520
rect 26635 2450 26650 2490
rect 26690 2450 26705 2490
rect 26635 2435 26705 2450
rect 27115 2490 27185 2520
rect 27115 2450 27130 2490
rect 27170 2450 27185 2490
rect 27115 2435 27185 2450
rect 28315 2490 28385 2520
rect 28315 2450 28330 2490
rect 28370 2450 28385 2490
rect 28315 2435 28385 2450
rect 30390 2490 30460 2520
rect 30390 2450 30405 2490
rect 30445 2450 30460 2490
rect 30390 2435 30460 2450
rect 31590 2490 31660 2520
rect 31590 2450 31605 2490
rect 31645 2450 31660 2490
rect 31590 2435 31660 2450
rect 32070 2490 32140 2520
rect 32070 2450 32085 2490
rect 32125 2450 32140 2490
rect 32070 2435 32140 2450
rect 33270 2490 33340 2520
rect 33270 2450 33285 2490
rect 33325 2450 33340 2490
rect 33270 2435 33340 2450
rect 35345 2490 35415 2520
rect 35345 2450 35360 2490
rect 35400 2450 35415 2490
rect 35345 2435 35415 2450
rect 36545 2490 36615 2520
rect 36545 2450 36560 2490
rect 36600 2450 36615 2490
rect 36545 2435 36615 2450
rect 37025 2490 37095 2520
rect 37025 2450 37040 2490
rect 37080 2450 37095 2490
rect 37025 2435 37095 2450
rect 38225 2490 38295 2520
rect 38225 2450 38240 2490
rect 38280 2450 38295 2490
rect 38225 2435 38295 2450
rect 40300 2490 40370 2520
rect 40300 2450 40315 2490
rect 40355 2450 40370 2490
rect 40300 2435 40370 2450
rect 41500 2490 41570 2520
rect 41500 2450 41515 2490
rect 41555 2450 41570 2490
rect 41500 2435 41570 2450
rect 41980 2490 42050 2520
rect 41980 2450 41995 2490
rect 42035 2450 42050 2490
rect 41980 2435 42050 2450
rect 43180 2490 43250 2520
rect 43180 2450 43195 2490
rect 43235 2450 43250 2490
rect 43180 2435 43250 2450
rect 45255 2490 45325 2520
rect 45255 2450 45270 2490
rect 45310 2450 45325 2490
rect 45255 2435 45325 2450
rect 46455 2490 46525 2520
rect 46455 2450 46470 2490
rect 46510 2450 46525 2490
rect 46455 2435 46525 2450
rect 46935 2490 47005 2520
rect 46935 2450 46950 2490
rect 46990 2450 47005 2490
rect 46935 2435 47005 2450
rect 48135 2490 48205 2520
rect 48135 2450 48150 2490
rect 48190 2450 48205 2490
rect 48135 2435 48205 2450
rect 50210 2490 50280 2520
rect 50210 2450 50225 2490
rect 50265 2450 50280 2490
rect 50210 2435 50280 2450
rect 51410 2490 51480 2520
rect 51410 2450 51425 2490
rect 51465 2450 51480 2490
rect 51410 2435 51480 2450
rect 51890 2490 51960 2520
rect 51890 2450 51905 2490
rect 51945 2450 51960 2490
rect 51890 2435 51960 2450
rect 53090 2490 53160 2520
rect 53090 2450 53105 2490
rect 53145 2450 53160 2490
rect 53090 2435 53160 2450
rect 55165 2490 55235 2520
rect 55165 2450 55180 2490
rect 55220 2450 55235 2490
rect 55165 2435 55235 2450
rect 56365 2490 56435 2520
rect 56365 2450 56380 2490
rect 56420 2450 56435 2490
rect 56365 2435 56435 2450
rect 56845 2490 56915 2520
rect 56845 2450 56860 2490
rect 56900 2450 56915 2490
rect 56845 2435 56915 2450
rect 58045 2490 58115 2520
rect 58045 2450 58060 2490
rect 58100 2450 58115 2490
rect 58045 2435 58115 2450
rect 60120 2490 60190 2520
rect 60120 2450 60135 2490
rect 60175 2450 60190 2490
rect 60120 2435 60190 2450
rect 61320 2490 61390 2520
rect 61320 2450 61335 2490
rect 61375 2450 61390 2490
rect 61320 2435 61390 2450
rect 61800 2490 61870 2520
rect 61800 2450 61815 2490
rect 61855 2450 61870 2490
rect 61800 2435 61870 2450
rect 63000 2490 63070 2520
rect 63000 2450 63015 2490
rect 63055 2450 63070 2490
rect 63000 2435 63070 2450
rect 65075 2490 65145 2520
rect 65075 2450 65090 2490
rect 65130 2450 65145 2490
rect 65075 2435 65145 2450
rect 66275 2490 66345 2520
rect 66275 2450 66290 2490
rect 66330 2450 66345 2490
rect 66275 2435 66345 2450
rect 66755 2490 66825 2520
rect 66755 2450 66770 2490
rect 66810 2450 66825 2490
rect 66755 2435 66825 2450
rect 67955 2490 68025 2520
rect 67955 2450 67970 2490
rect 68010 2450 68025 2490
rect 67955 2435 68025 2450
rect 70030 2490 70100 2520
rect 70030 2450 70045 2490
rect 70085 2450 70100 2490
rect 70030 2435 70100 2450
rect 71230 2490 71300 2520
rect 71230 2450 71245 2490
rect 71285 2450 71300 2490
rect 71230 2435 71300 2450
rect 71710 2490 71780 2520
rect 71710 2450 71725 2490
rect 71765 2450 71780 2490
rect 71710 2435 71780 2450
rect 72910 2490 72980 2520
rect 72910 2450 72925 2490
rect 72965 2450 72980 2490
rect 72910 2435 72980 2450
rect 74985 2490 75055 2520
rect 74985 2450 75000 2490
rect 75040 2450 75055 2490
rect 74985 2435 75055 2450
rect 76185 2490 76255 2520
rect 76185 2450 76200 2490
rect 76240 2450 76255 2490
rect 76185 2435 76255 2450
rect 76665 2490 76735 2520
rect 76665 2450 76680 2490
rect 76720 2450 76735 2490
rect 76665 2435 76735 2450
rect 77865 2490 77935 2520
rect 77865 2450 77880 2490
rect 77920 2450 77935 2490
rect 77865 2435 77935 2450
rect -345 2405 -280 2420
rect -345 2370 -330 2405
rect -295 2385 -280 2405
rect -295 2370 0 2385
rect -345 2355 0 2370
rect 4295 2355 4955 2385
rect 9250 2355 9910 2385
rect 14205 2355 14865 2385
rect 19160 2355 19820 2385
rect 24115 2355 24775 2385
rect 29070 2355 29730 2385
rect 34025 2355 34685 2385
rect 38980 2355 39640 2385
rect 43935 2355 44595 2385
rect 48890 2355 49550 2385
rect 53845 2355 54505 2385
rect 58800 2355 59460 2385
rect 63755 2355 64415 2385
rect 68710 2355 69370 2385
rect 73665 2355 74325 2385
rect 8690 2250 8775 2265
rect 8690 2210 8705 2250
rect 8745 2210 8775 2250
rect 8690 2195 8775 2210
rect 10355 2250 10440 2265
rect 10355 2210 10385 2250
rect 10425 2210 10440 2250
rect 10355 2195 10440 2210
rect 13645 2250 13730 2265
rect 13645 2210 13660 2250
rect 13700 2210 13730 2250
rect 13645 2195 13730 2210
rect 15310 2250 15395 2265
rect 15310 2210 15340 2250
rect 15380 2210 15395 2250
rect 15310 2195 15395 2210
rect 18600 2250 18685 2265
rect 18600 2210 18615 2250
rect 18655 2210 18685 2250
rect 18600 2195 18685 2210
rect 20265 2250 20350 2265
rect 20265 2210 20295 2250
rect 20335 2210 20350 2250
rect 20265 2195 20350 2210
rect 23555 2250 23640 2265
rect 23555 2210 23570 2250
rect 23610 2210 23640 2250
rect 23555 2195 23640 2210
rect 25220 2250 25305 2265
rect 25220 2210 25250 2250
rect 25290 2210 25305 2250
rect 25220 2195 25305 2210
rect 28510 2250 28595 2265
rect 28510 2210 28525 2250
rect 28565 2210 28595 2250
rect 28510 2195 28595 2210
rect 30175 2250 30260 2265
rect 30175 2210 30205 2250
rect 30245 2210 30260 2250
rect 30175 2195 30260 2210
rect 33465 2250 33550 2265
rect 33465 2210 33480 2250
rect 33520 2210 33550 2250
rect 33465 2195 33550 2210
rect 35130 2250 35215 2265
rect 35130 2210 35160 2250
rect 35200 2210 35215 2250
rect 35130 2195 35215 2210
rect 38420 2250 38505 2265
rect 38420 2210 38435 2250
rect 38475 2210 38505 2250
rect 38420 2195 38505 2210
rect 40085 2250 40170 2265
rect 40085 2210 40115 2250
rect 40155 2210 40170 2250
rect 40085 2195 40170 2210
rect 43375 2250 43460 2265
rect 43375 2210 43390 2250
rect 43430 2210 43460 2250
rect 43375 2195 43460 2210
rect 45040 2250 45125 2265
rect 45040 2210 45070 2250
rect 45110 2210 45125 2250
rect 45040 2195 45125 2210
rect 48330 2250 48415 2265
rect 48330 2210 48345 2250
rect 48385 2210 48415 2250
rect 48330 2195 48415 2210
rect 49995 2250 50080 2265
rect 49995 2210 50025 2250
rect 50065 2210 50080 2250
rect 49995 2195 50080 2210
rect 53285 2250 53370 2265
rect 53285 2210 53300 2250
rect 53340 2210 53370 2250
rect 53285 2195 53370 2210
rect 54950 2250 55035 2265
rect 54950 2210 54980 2250
rect 55020 2210 55035 2250
rect 54950 2195 55035 2210
rect 58240 2250 58325 2265
rect 58240 2210 58255 2250
rect 58295 2210 58325 2250
rect 58240 2195 58325 2210
rect 59905 2250 59990 2265
rect 59905 2210 59935 2250
rect 59975 2210 59990 2250
rect 59905 2195 59990 2210
rect 63195 2250 63280 2265
rect 63195 2210 63210 2250
rect 63250 2210 63280 2250
rect 63195 2195 63280 2210
rect 64860 2250 64945 2265
rect 64860 2210 64890 2250
rect 64930 2210 64945 2250
rect 64860 2195 64945 2210
rect 68150 2250 68235 2265
rect 68150 2210 68165 2250
rect 68205 2210 68235 2250
rect 68150 2195 68235 2210
rect 69815 2250 69900 2265
rect 69815 2210 69845 2250
rect 69885 2210 69900 2250
rect 69815 2195 69900 2210
rect 73105 2250 73190 2265
rect 73105 2210 73120 2250
rect 73160 2210 73190 2250
rect 73105 2195 73190 2210
rect 74770 2250 74855 2265
rect 74770 2210 74800 2250
rect 74840 2210 74855 2250
rect 74770 2195 74855 2210
rect 8690 330 8775 345
rect 8690 290 8705 330
rect 8745 290 8775 330
rect 8690 275 8775 290
rect 10355 330 10440 345
rect 10355 290 10385 330
rect 10425 290 10440 330
rect 10355 275 10440 290
rect 13645 330 13730 345
rect 13645 290 13660 330
rect 13700 290 13730 330
rect 13645 275 13730 290
rect 15310 330 15395 345
rect 15310 290 15340 330
rect 15380 290 15395 330
rect 15310 275 15395 290
rect 18600 330 18685 345
rect 18600 290 18615 330
rect 18655 290 18685 330
rect 18600 275 18685 290
rect 20265 330 20350 345
rect 20265 290 20295 330
rect 20335 290 20350 330
rect 20265 275 20350 290
rect 23555 330 23640 345
rect 23555 290 23570 330
rect 23610 290 23640 330
rect 23555 275 23640 290
rect 25220 330 25305 345
rect 25220 290 25250 330
rect 25290 290 25305 330
rect 25220 275 25305 290
rect 28510 330 28595 345
rect 28510 290 28525 330
rect 28565 290 28595 330
rect 28510 275 28595 290
rect 30175 330 30260 345
rect 30175 290 30205 330
rect 30245 290 30260 330
rect 30175 275 30260 290
rect 33465 330 33550 345
rect 33465 290 33480 330
rect 33520 290 33550 330
rect 33465 275 33550 290
rect 35130 330 35215 345
rect 35130 290 35160 330
rect 35200 290 35215 330
rect 35130 275 35215 290
rect 38420 330 38505 345
rect 38420 290 38435 330
rect 38475 290 38505 330
rect 38420 275 38505 290
rect 40085 330 40170 345
rect 40085 290 40115 330
rect 40155 290 40170 330
rect 40085 275 40170 290
rect 43375 330 43460 345
rect 43375 290 43390 330
rect 43430 290 43460 330
rect 43375 275 43460 290
rect 45040 330 45125 345
rect 45040 290 45070 330
rect 45110 290 45125 330
rect 45040 275 45125 290
rect 48330 330 48415 345
rect 48330 290 48345 330
rect 48385 290 48415 330
rect 48330 275 48415 290
rect 49995 330 50080 345
rect 49995 290 50025 330
rect 50065 290 50080 330
rect 49995 275 50080 290
rect 53285 330 53370 345
rect 53285 290 53300 330
rect 53340 290 53370 330
rect 53285 275 53370 290
rect 54950 330 55035 345
rect 54950 290 54980 330
rect 55020 290 55035 330
rect 54950 275 55035 290
rect 58240 330 58325 345
rect 58240 290 58255 330
rect 58295 290 58325 330
rect 58240 275 58325 290
rect 59905 330 59990 345
rect 59905 290 59935 330
rect 59975 290 59990 330
rect 59905 275 59990 290
rect 63195 330 63280 345
rect 63195 290 63210 330
rect 63250 290 63280 330
rect 63195 275 63280 290
rect 64860 330 64945 345
rect 64860 290 64890 330
rect 64930 290 64945 330
rect 64860 275 64945 290
rect 68150 330 68235 345
rect 68150 290 68165 330
rect 68205 290 68235 330
rect 68150 275 68235 290
rect 69815 330 69900 345
rect 69815 290 69845 330
rect 69885 290 69900 330
rect 69815 275 69900 290
rect 73105 330 73190 345
rect 73105 290 73120 330
rect 73160 290 73190 330
rect 73105 275 73190 290
rect 74770 330 74855 345
rect 74770 290 74800 330
rect 74840 290 74855 330
rect 74770 275 74855 290
rect 15 185 80 200
rect 15 150 30 185
rect 65 150 80 185
rect 15 135 80 150
rect 4365 135 4970 165
rect 9320 135 9925 165
rect 14275 135 14880 165
rect 19230 135 19835 165
rect 24185 135 24790 165
rect 29140 135 29745 165
rect 34095 135 34700 165
rect 39050 135 39655 165
rect 44005 135 44610 165
rect 48960 135 49565 165
rect 53915 135 54520 165
rect 58870 135 59475 165
rect 63825 135 64430 165
rect 68780 135 69385 165
rect 73735 135 74340 165
<< via1 >>
rect -330 11595 -295 11630
rect 30 9375 65 9410
rect -330 8520 -295 8555
rect 30 6300 65 6335
rect -330 5445 -295 5480
rect 30 3225 65 3260
rect -330 2370 -295 2405
rect 30 150 65 185
<< metal2 >>
rect -345 11630 -280 11645
rect -345 11595 -330 11630
rect -295 11595 -280 11630
rect -345 8555 -280 11595
rect -345 8520 -330 8555
rect -295 8520 -280 8555
rect -345 5480 -280 8520
rect -345 5445 -330 5480
rect -295 5445 -280 5480
rect -345 2405 -280 5445
rect -345 2370 -330 2405
rect -295 2370 -280 2405
rect -345 2355 -280 2370
rect 15 9410 80 9425
rect 15 9375 30 9410
rect 65 9375 80 9410
rect 15 6335 80 9375
rect 15 6300 30 6335
rect 65 6300 80 6335
rect 15 3260 80 6300
rect 15 3225 30 3260
rect 65 3225 80 3260
rect 15 1310 80 3225
rect -345 1255 80 1310
rect 15 185 80 1255
rect 15 150 30 185
rect 65 150 80 185
rect 15 135 80 150
use nmos_final_middle  nmos_final_middle_0
array 0 15 4955 0 3 3075
timestamp 1641483920
transform 1 0 1065 0 1 -9985
box -1065 9960 3300 12505
<< labels >>
rlabel metal1 -345 11985 -345 11985 7 G
port 1 w
rlabel metal2 -345 11610 -345 11610 7 D
port 2 w
rlabel metal2 -345 1280 -345 1280 7 S
port 3 w
rlabel locali -345 1740 -345 1740 7 B
port 4 w
<< end >>
