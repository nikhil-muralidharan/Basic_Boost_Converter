magic
tech sky130A
timestamp 1660237895
<< nwell >>
rect 1130 220 1900 385
rect 180 -440 1035 -220
<< pmoslvt >>
rect 335 -385 370 -285
rect 510 -385 545 -285
rect 595 -385 630 -285
<< nmoslvt >>
rect 185 -590 200 -490
rect 335 -590 350 -490
rect 510 -590 525 -490
rect 660 -590 675 -490
<< ndiff >>
rect 135 -505 185 -490
rect 135 -575 150 -505
rect 170 -575 185 -505
rect 135 -590 185 -575
rect 200 -505 250 -490
rect 200 -575 215 -505
rect 235 -575 250 -505
rect 200 -590 250 -575
rect 285 -505 335 -490
rect 285 -575 300 -505
rect 320 -575 335 -505
rect 285 -590 335 -575
rect 350 -505 400 -490
rect 350 -575 365 -505
rect 385 -575 400 -505
rect 350 -590 400 -575
rect 460 -505 510 -490
rect 460 -575 475 -505
rect 495 -575 510 -505
rect 460 -590 510 -575
rect 525 -505 575 -490
rect 525 -575 540 -505
rect 560 -575 575 -505
rect 525 -590 575 -575
rect 610 -505 660 -490
rect 610 -575 625 -505
rect 645 -575 660 -505
rect 610 -590 660 -575
rect 675 -505 725 -490
rect 675 -575 690 -505
rect 710 -575 725 -505
rect 675 -590 725 -575
<< pdiff >>
rect 285 -300 335 -285
rect 285 -370 300 -300
rect 320 -370 335 -300
rect 285 -385 335 -370
rect 370 -300 420 -285
rect 370 -370 385 -300
rect 405 -370 420 -300
rect 370 -385 420 -370
rect 460 -300 510 -285
rect 460 -370 475 -300
rect 495 -370 510 -300
rect 460 -385 510 -370
rect 545 -300 595 -285
rect 545 -370 560 -300
rect 580 -370 595 -300
rect 545 -385 595 -370
rect 630 -300 680 -285
rect 630 -370 645 -300
rect 665 -370 680 -300
rect 630 -385 680 -370
<< ndiffc >>
rect 150 -575 170 -505
rect 215 -575 235 -505
rect 300 -575 320 -505
rect 365 -575 385 -505
rect 475 -575 495 -505
rect 540 -575 560 -505
rect 625 -575 645 -505
rect 690 -575 710 -505
<< pdiffc >>
rect 300 -370 320 -300
rect 385 -370 405 -300
rect 475 -370 495 -300
rect 560 -370 580 -300
rect 645 -370 665 -300
<< psubdiff >>
rect 15 -505 65 -490
rect 15 -575 30 -505
rect 50 -575 65 -505
rect 15 -590 65 -575
<< nsubdiff >>
rect 200 -300 250 -285
rect 200 -370 215 -300
rect 235 -370 250 -300
rect 200 -385 250 -370
<< psubdiffcont >>
rect 30 -575 50 -505
<< nsubdiffcont >>
rect 215 -370 235 -300
<< poly >>
rect 335 -240 375 -230
rect 335 -260 345 -240
rect 365 -260 375 -240
rect 335 -270 375 -260
rect 505 -240 545 -230
rect 505 -260 515 -240
rect 535 -260 545 -240
rect 505 -270 545 -260
rect 335 -285 370 -270
rect 510 -285 545 -270
rect 595 -285 630 -270
rect 335 -400 370 -385
rect 510 -400 545 -385
rect 595 -400 630 -385
rect 335 -410 375 -400
rect 335 -430 345 -410
rect 365 -430 375 -410
rect 335 -440 375 -430
rect 590 -410 630 -400
rect 590 -430 600 -410
rect 620 -430 630 -410
rect 590 -440 630 -430
rect 185 -490 200 -475
rect 335 -490 350 -475
rect 510 -490 525 -475
rect 660 -490 675 -475
rect 185 -605 200 -590
rect 335 -605 350 -590
rect 510 -605 525 -590
rect 660 -605 675 -590
rect 185 -615 225 -605
rect 185 -635 195 -615
rect 215 -635 225 -615
rect 185 -645 225 -635
rect 335 -615 375 -605
rect 335 -635 345 -615
rect 365 -635 375 -615
rect 335 -645 375 -635
rect 510 -615 550 -605
rect 510 -635 520 -615
rect 540 -635 550 -615
rect 510 -645 550 -635
rect 660 -615 700 -605
rect 660 -635 670 -615
rect 690 -635 700 -615
rect 660 -645 700 -635
<< polycont >>
rect 345 -260 365 -240
rect 515 -260 535 -240
rect 345 -430 365 -410
rect 600 -430 620 -410
rect 195 -635 215 -615
rect 345 -635 365 -615
rect 520 -635 540 -615
rect 670 -635 690 -615
<< locali >>
rect 520 20 670 40
rect 1135 20 1270 40
rect 400 -25 420 10
rect 825 -25 845 10
rect 400 -45 845 -25
rect 1450 -70 1470 10
rect 1055 -90 1470 -70
rect 5 -170 590 -150
rect 5 -220 310 -200
rect 290 -290 310 -220
rect 335 -240 375 -230
rect 505 -240 545 -230
rect 335 -260 345 -240
rect 365 -260 515 -240
rect 535 -260 545 -240
rect 335 -270 375 -260
rect 505 -270 545 -260
rect 570 -290 590 -170
rect 205 -300 245 -290
rect 205 -370 215 -300
rect 235 -370 245 -300
rect 205 -380 245 -370
rect 290 -300 330 -290
rect 290 -370 300 -300
rect 320 -370 330 -300
rect 290 -380 330 -370
rect 375 -300 415 -290
rect 375 -370 385 -300
rect 405 -370 415 -300
rect 375 -380 415 -370
rect 465 -300 505 -290
rect 465 -370 475 -300
rect 495 -370 505 -300
rect 465 -380 505 -370
rect 550 -300 590 -290
rect 550 -370 560 -300
rect 580 -370 590 -300
rect 550 -380 590 -370
rect 635 -300 675 -290
rect 635 -370 645 -300
rect 665 -370 675 -300
rect 635 -380 675 -370
rect 300 -400 320 -380
rect 300 -410 375 -400
rect 300 -430 345 -410
rect 365 -430 375 -410
rect 300 -440 375 -430
rect 475 -410 495 -380
rect 655 -400 675 -380
rect 590 -410 630 -400
rect 475 -430 600 -410
rect 620 -430 630 -410
rect 655 -420 710 -400
rect 300 -495 320 -440
rect 475 -495 495 -430
rect 590 -440 630 -430
rect 690 -495 710 -420
rect 20 -505 60 -495
rect 20 -575 30 -505
rect 50 -575 60 -505
rect 20 -585 60 -575
rect 140 -505 180 -495
rect 140 -575 150 -505
rect 170 -575 180 -505
rect 140 -585 180 -575
rect 205 -505 245 -495
rect 205 -575 215 -505
rect 235 -575 245 -505
rect 205 -585 245 -575
rect 290 -505 330 -495
rect 290 -575 300 -505
rect 320 -575 330 -505
rect 290 -585 330 -575
rect 355 -505 395 -495
rect 355 -575 365 -505
rect 385 -575 395 -505
rect 355 -585 395 -575
rect 465 -505 505 -495
rect 465 -575 475 -505
rect 495 -575 505 -505
rect 465 -585 505 -575
rect 530 -505 570 -495
rect 530 -575 540 -505
rect 560 -575 570 -505
rect 530 -585 570 -575
rect 615 -505 655 -495
rect 615 -575 625 -505
rect 645 -575 655 -505
rect 615 -585 655 -575
rect 680 -505 720 -495
rect 680 -575 690 -505
rect 710 -575 720 -505
rect 680 -585 720 -575
rect 215 -605 235 -585
rect 1055 -605 1075 -90
rect 185 -615 235 -605
rect 335 -615 375 -605
rect 510 -615 550 -605
rect 660 -615 700 -605
rect 185 -635 195 -615
rect 215 -635 345 -615
rect 365 -635 520 -615
rect 540 -635 670 -615
rect 690 -635 700 -615
rect 1035 -625 1075 -605
rect 185 -645 225 -635
rect 335 -645 375 -635
rect 510 -645 550 -635
rect 660 -645 700 -635
<< viali >>
rect 215 -370 235 -300
rect 30 -575 50 -505
rect 150 -575 170 -505
rect 365 -575 385 -505
rect 540 -575 560 -505
rect 625 -575 645 -505
<< metal1 >>
rect 195 -300 255 -290
rect 195 -370 215 -300
rect 235 -370 255 -300
rect 195 -380 255 -370
rect 185 -495 200 -490
rect 335 -495 350 -490
rect 510 -495 525 -490
rect 660 -495 675 -490
rect 5 -505 775 -495
rect 5 -575 30 -505
rect 50 -575 150 -505
rect 170 -575 365 -505
rect 385 -575 540 -505
rect 560 -575 625 -505
rect 645 -575 775 -505
rect 5 -585 775 -575
rect 185 -590 200 -585
rect 335 -590 350 -585
rect 510 -590 525 -585
rect 660 -590 675 -585
use inverter_lvt_zcd  inverter_lvt_zcd_0
timestamp 1658301810
transform 1 0 185 0 1 80
box -185 -80 75 300
use inverter_lvt_zcd  inverter_lvt_zcd_1
timestamp 1658301810
transform 1 0 445 0 1 80
box -185 -80 75 300
use inverter_lvt_zcd  inverter_lvt_zcd_2
timestamp 1658301810
transform 1 0 960 0 1 -565
box -185 -80 75 300
use or_lvt_zcd  or_lvt_zcd_0
timestamp 1659680843
transform 1 0 725 0 1 105
box -205 -105 410 280
use sr_latch_lvt_zcd  sr_latch_lvt_zcd_0
timestamp 1660234770
transform 1 0 1410 0 1 130
box -280 -130 500 240
<< end >>
