magic
tech sky130A
timestamp 1660757217
<< nwell >>
rect -185 140 75 300
<< pmoslvt >>
rect -30 170 5 270
<< nmoslvt >>
rect -30 -300 -15 -200
<< ndiff >>
rect -80 -215 -30 -200
rect -80 -285 -65 -215
rect -45 -285 -30 -215
rect -80 -300 -30 -285
rect -15 -215 35 -200
rect -15 -285 0 -215
rect 20 -285 35 -215
rect -15 -300 35 -285
<< pdiff >>
rect -80 255 -30 270
rect -80 185 -65 255
rect -45 185 -30 255
rect -80 170 -30 185
rect 5 255 55 270
rect 5 185 20 255
rect 40 185 55 255
rect 5 170 55 185
<< ndiffc >>
rect -65 -285 -45 -215
rect 0 -285 20 -215
<< pdiffc >>
rect -65 185 -45 255
rect 20 185 40 255
<< psubdiff >>
rect -165 -215 -115 -200
rect -165 -285 -150 -215
rect -130 -285 -115 -215
rect -165 -300 -115 -285
<< nsubdiff >>
rect -165 255 -115 270
rect -165 185 -150 255
rect -130 185 -115 255
rect -165 170 -115 185
<< psubdiffcont >>
rect -150 -285 -130 -215
<< nsubdiffcont >>
rect -150 185 -130 255
<< poly >>
rect -30 270 5 285
rect -30 155 5 170
rect -30 80 -15 155
rect -55 70 -15 80
rect -55 50 -45 70
rect -25 50 -15 70
rect -55 40 -15 50
rect -55 -155 -15 -145
rect -55 -175 -45 -155
rect -25 -175 -15 -155
rect -55 -185 -15 -175
rect -30 -200 -15 -185
rect -30 -315 -15 -300
rect -55 -325 -15 -315
rect -55 -345 -45 -325
rect -25 -345 -15 -325
rect -55 -355 -15 -345
<< polycont >>
rect -45 50 -25 70
rect -45 -175 -25 -155
rect -45 -345 -25 -325
<< locali >>
rect -160 255 -120 265
rect -160 185 -150 255
rect -130 185 -120 255
rect -160 175 -120 185
rect -75 255 -35 265
rect -75 185 -65 255
rect -45 185 -35 255
rect -75 175 -35 185
rect 10 255 50 265
rect 10 185 20 255
rect 40 185 50 255
rect 10 175 50 185
rect -55 70 -15 80
rect -55 50 -45 70
rect -25 50 -15 70
rect -55 40 -15 50
rect -45 -145 -25 40
rect -55 -155 -15 -145
rect -55 -175 -45 -155
rect -25 -175 -15 -155
rect -55 -185 -15 -175
rect 10 -205 30 175
rect -160 -215 -120 -205
rect -160 -285 -150 -215
rect -130 -285 -120 -215
rect -160 -295 -120 -285
rect -75 -215 -35 -205
rect -75 -285 -65 -215
rect -45 -285 -35 -215
rect -75 -295 -35 -285
rect -10 -215 30 -205
rect -10 -285 0 -215
rect 20 -285 30 -215
rect -10 -295 30 -285
rect 10 -315 30 -295
rect -185 -325 -15 -315
rect -185 -335 -45 -325
rect -55 -345 -45 -335
rect -25 -345 -15 -325
rect 10 -335 75 -315
rect -55 -355 -15 -345
<< viali >>
rect -150 185 -130 255
rect -65 185 -45 255
rect -150 -285 -130 -215
rect -65 -285 -45 -215
<< metal1 >>
rect -185 255 75 265
rect -185 185 -150 255
rect -130 185 -65 255
rect -45 185 75 255
rect -185 175 75 185
rect -185 -215 75 -205
rect -185 -285 -150 -215
rect -130 -285 -65 -215
rect -45 -285 75 -215
rect -185 -295 75 -285
<< labels >>
rlabel metal1 -185 220 -185 220 7 VP
port 3 w
rlabel metal1 -185 -250 -185 -250 7 VN
port 4 w
rlabel locali -185 -325 -185 -325 7 in
port 1 w
rlabel locali 75 -320 75 -320 3 out
port 2 e
<< end >>
