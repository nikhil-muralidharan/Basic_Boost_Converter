magic
tech sky130A
timestamp 1660758955
<< nwell >>
rect -160 220 490 380
<< pmoslvt >>
rect 0 250 35 350
rect 165 250 200 350
rect 330 250 365 350
<< nmoslvt >>
rect 55 -220 70 -120
rect 120 -220 135 -120
rect 265 -220 280 -120
<< ndiff >>
rect 5 -135 55 -120
rect 5 -205 20 -135
rect 40 -205 55 -135
rect 5 -220 55 -205
rect 70 -135 120 -120
rect 70 -205 85 -135
rect 105 -205 120 -135
rect 70 -220 120 -205
rect 135 -135 185 -120
rect 135 -205 150 -135
rect 170 -205 185 -135
rect 135 -220 185 -205
rect 215 -135 265 -120
rect 215 -205 230 -135
rect 250 -205 265 -135
rect 215 -220 265 -205
rect 280 -135 330 -120
rect 280 -205 295 -135
rect 315 -205 330 -135
rect 280 -220 330 -205
<< pdiff >>
rect -50 335 0 350
rect -50 265 -35 335
rect -15 265 0 335
rect -50 250 0 265
rect 35 335 85 350
rect 35 265 50 335
rect 70 265 85 335
rect 35 250 85 265
rect 115 335 165 350
rect 115 265 130 335
rect 150 265 165 335
rect 115 250 165 265
rect 200 335 250 350
rect 200 265 215 335
rect 235 265 250 335
rect 200 250 250 265
rect 280 335 330 350
rect 280 265 295 335
rect 315 265 330 335
rect 280 250 330 265
rect 365 335 415 350
rect 365 265 380 335
rect 400 265 415 335
rect 365 250 415 265
<< ndiffc >>
rect 20 -205 40 -135
rect 85 -205 105 -135
rect 150 -205 170 -135
rect 230 -205 250 -135
rect 295 -205 315 -135
<< pdiffc >>
rect -35 265 -15 335
rect 50 265 70 335
rect 130 265 150 335
rect 215 265 235 335
rect 295 265 315 335
rect 380 265 400 335
<< psubdiff >>
rect -75 -130 -25 -120
rect -75 -205 -60 -130
rect -40 -205 -25 -130
rect -75 -220 -25 -205
<< nsubdiff >>
rect -130 340 -80 350
rect -130 265 -115 340
rect -95 265 -80 340
rect -130 250 -80 265
<< psubdiffcont >>
rect -60 -205 -40 -130
<< nsubdiffcont >>
rect -115 265 -95 340
<< poly >>
rect 0 395 40 405
rect 0 375 10 395
rect 30 375 40 395
rect 0 365 40 375
rect 165 395 205 405
rect 165 375 175 395
rect 195 375 205 395
rect 165 365 205 375
rect 0 350 35 365
rect 165 350 200 365
rect 330 350 365 365
rect 0 240 35 250
rect 165 240 200 250
rect 330 240 365 250
rect 0 225 70 240
rect 55 175 70 225
rect 120 225 200 240
rect 265 225 365 240
rect 120 175 135 225
rect 265 215 280 225
rect 240 205 280 215
rect 240 185 250 205
rect 270 185 280 205
rect 240 175 280 185
rect 35 165 75 175
rect 35 145 45 165
rect 65 145 75 165
rect 35 135 75 145
rect 120 165 160 175
rect 120 145 130 165
rect 150 145 160 165
rect 120 135 160 145
rect 55 -70 95 -60
rect 55 -90 65 -70
rect 85 -90 95 -70
rect 55 -100 95 -90
rect 120 -70 160 -60
rect 120 -90 130 -70
rect 150 -90 160 -70
rect 120 -100 160 -90
rect 240 -70 280 -60
rect 240 -90 250 -70
rect 270 -90 280 -70
rect 240 -100 280 -90
rect 55 -120 70 -100
rect 120 -120 135 -100
rect 265 -120 280 -100
rect 55 -235 70 -220
rect 30 -245 70 -235
rect 30 -265 40 -245
rect 60 -265 70 -245
rect 30 -275 70 -265
rect 120 -235 135 -220
rect 265 -235 280 -220
rect 120 -245 160 -235
rect 120 -265 130 -245
rect 150 -265 160 -245
rect 120 -275 160 -265
<< polycont >>
rect 10 375 30 395
rect 175 375 195 395
rect 250 185 270 205
rect 45 145 65 165
rect 130 145 150 165
rect 65 -90 85 -70
rect 130 -90 150 -70
rect 250 -90 270 -70
rect 40 -265 60 -245
rect 130 -265 150 -245
<< locali >>
rect 0 395 40 405
rect 0 375 10 395
rect 30 375 40 395
rect 0 365 40 375
rect 165 395 205 405
rect 165 375 175 395
rect 195 375 205 395
rect 165 365 205 375
rect -125 340 -85 345
rect -125 265 -115 340
rect -95 265 -85 340
rect -125 255 -85 265
rect -45 335 -5 345
rect -45 265 -35 335
rect -15 265 -5 335
rect -45 255 -5 265
rect 40 335 80 345
rect 40 265 50 335
rect 70 265 80 335
rect 40 255 80 265
rect 120 335 160 345
rect 120 265 130 335
rect 150 265 160 335
rect 120 255 160 265
rect 205 335 245 345
rect 205 265 215 335
rect 235 265 245 335
rect 205 255 245 265
rect 285 335 325 345
rect 285 265 295 335
rect 315 265 325 335
rect 285 255 325 265
rect 370 335 410 345
rect 370 265 380 335
rect 400 265 410 335
rect 370 255 410 265
rect -35 215 -15 255
rect 130 215 150 255
rect -35 205 280 215
rect -35 195 250 205
rect -35 -75 -15 195
rect 240 185 250 195
rect 270 185 280 205
rect 240 175 280 185
rect 300 205 320 255
rect 300 185 435 205
rect 35 165 75 175
rect 35 145 45 165
rect 65 145 75 165
rect 35 135 75 145
rect 120 165 160 175
rect 120 145 130 165
rect 150 145 160 165
rect 120 135 160 145
rect 55 -60 75 135
rect 130 -60 150 135
rect 250 -60 270 175
rect 55 -70 95 -60
rect -35 -95 30 -75
rect 10 -125 30 -95
rect 55 -90 65 -70
rect 85 -90 95 -70
rect 55 -100 95 -90
rect 120 -70 160 -60
rect 120 -90 130 -70
rect 150 -90 160 -70
rect 120 -100 160 -90
rect 240 -70 280 -60
rect 240 -90 250 -70
rect 270 -90 280 -70
rect 240 -100 280 -90
rect 300 -125 320 185
rect -70 -130 -30 -125
rect -70 -205 -60 -130
rect -40 -205 -30 -130
rect -70 -215 -30 -205
rect 10 -135 50 -125
rect 10 -205 20 -135
rect 40 -205 50 -135
rect 10 -215 50 -205
rect 75 -135 115 -125
rect 75 -205 85 -135
rect 105 -205 115 -135
rect 75 -215 115 -205
rect 140 -135 180 -125
rect 140 -205 150 -135
rect 170 -205 180 -135
rect 140 -215 180 -205
rect 220 -135 260 -125
rect 220 -205 230 -135
rect 250 -205 260 -135
rect 220 -215 260 -205
rect 285 -135 325 -125
rect 285 -205 295 -135
rect 315 -205 325 -135
rect 285 -215 325 -205
rect 415 -235 435 185
rect 30 -245 70 -235
rect 30 -265 40 -245
rect 60 -265 70 -245
rect 30 -275 70 -265
rect 120 -245 160 -235
rect 120 -265 130 -245
rect 150 -265 160 -245
rect 415 -255 500 -235
rect 120 -275 160 -265
<< viali >>
rect -115 265 -95 340
rect 50 265 70 335
rect 215 265 235 335
rect 380 265 400 335
rect -60 -205 -40 -130
rect 150 -205 170 -135
rect 230 -205 250 -135
<< metal1 >>
rect -160 340 490 345
rect -160 265 -115 340
rect -95 335 490 340
rect -95 265 50 335
rect 70 265 215 335
rect 235 265 380 335
rect 400 265 490 335
rect -160 255 490 265
rect -160 -130 490 -125
rect -160 -205 -60 -130
rect -40 -135 490 -130
rect -40 -205 150 -135
rect 170 -205 230 -135
rect 250 -205 490 -135
rect -160 -215 490 -205
<< labels >>
rlabel locali 435 195 435 195 3 Y
port 5 e
rlabel metal1 -160 300 -160 300 7 VP
port 1 w
rlabel locali 20 405 20 405 1 A
port 3 n
rlabel locali 185 405 185 405 1 B
port 4 n
rlabel metal1 -160 -165 -160 -165 7 VN
port 2 w
<< end >>
