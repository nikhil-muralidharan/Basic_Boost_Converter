**.subckt Basic_Boost
C1 Vout GND 4.375u m=1
R1 Vout GND 6 m=1
L1 Vin net1 3.125u m=1
V1 Vin GND pwl 0 1 0.25ms 1 0.251ms 1.2 0.500ms 1.2 0.501ms 1.4
V2 Ndrive GND PULSE (0 1 0 0.01us 0.01us 0.85us 1.25us)
V3 Pdrive GND PULSE (0 1 0 0.01us 0.01us 0.85us 1.25us)
X1 Ndrive net1 GND powern
X2 Pdrive net1 Vout powerp
**** begin user architecture code
** manual skywater pdks install (with patches applied)
* .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt_mm

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt_mm




.tran 0.1ms 1ms
.save all
.option savecurrents

**** end user architecture code
**.ends

* expanding   symbol:  powern.sym # of pins=3
** sym_path: /home/nikhil/Desktop/Basic_Boost_Converter/Spice_Files/powern.sym
** sch_path: /home/nikhil/Desktop/Basic_Boost_Converter/Spice_Files/powern.sch
.subckt powern  NDRIVE VDDIN VSSOUT
X0 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X2 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X3 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X4 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X5 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X6 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X7 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X8 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X9 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X10 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X11 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X12 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X13 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X14 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X15 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X16 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X17 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X18 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X19 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X20 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X21 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X22 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X23 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X24 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X25 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X26 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X27 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X28 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X29 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X30 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X31 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X32 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X33 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X34 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X35 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X36 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X37 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X38 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X39 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X40 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X41 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X42 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X43 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X44 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X45 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X46 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X47 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X48 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X49 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X50 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X51 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X52 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X53 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X54 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X55 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X56 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X57 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X58 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X59 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X60 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X61 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X62 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X63 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X64 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X65 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X66 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X67 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X68 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X69 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X70 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X71 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X72 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X73 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X74 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X75 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X76 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X77 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X78 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X79 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X80 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X81 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X82 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X83 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X84 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X85 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X86 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X87 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X88 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X89 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X90 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X91 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X92 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X93 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X94 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X95 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X96 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X97 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X98 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X99 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X100 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X101 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X102 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X103 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X104 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X105 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X106 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X107 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X108 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X109 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X110 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X111 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X112 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X113 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X114 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X115 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X116 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X117 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X118 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X119 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X120 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X121 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X122 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X123 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X124 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X125 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X126 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X127 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X128 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X129 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X130 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X131 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X132 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X133 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X134 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X135 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X136 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X137 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X138 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X139 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X140 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X141 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X142 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X143 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X144 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X145 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X146 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X147 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X148 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X149 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X150 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X151 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X152 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X153 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X154 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X155 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X156 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X157 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X158 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X159 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X160 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X161 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X162 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X163 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X164 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X165 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X166 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X167 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X168 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X169 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X170 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X171 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X172 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X173 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X174 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X175 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X176 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X177 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X178 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X179 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X180 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X181 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X182 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X183 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X184 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X185 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X186 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X187 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X188 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X189 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X190 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X191 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X192 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X193 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X194 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X195 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X196 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X197 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X198 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X199 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X200 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X201 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X202 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X203 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X204 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X205 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X206 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X207 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X208 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X209 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X210 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X211 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X212 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X213 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X214 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X215 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X216 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X217 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X218 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X219 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X220 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X221 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X222 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X223 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X224 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X225 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X226 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X227 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X228 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X229 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X230 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X231 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X232 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X233 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X234 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X235 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X236 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X237 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X238 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X239 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X240 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X241 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X242 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X243 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X244 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X245 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X246 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X247 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X248 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X249 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X250 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X251 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X252 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X253 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X254 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X255 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X256 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X257 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X258 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X259 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X260 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X261 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X262 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X263 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X264 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X265 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X266 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X267 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X268 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X269 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X270 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X271 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X272 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X273 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X274 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X275 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X276 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X277 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X278 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X279 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X280 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X281 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X282 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X283 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X284 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X285 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X286 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X287 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X288 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X289 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X290 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X291 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X292 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X293 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X294 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X295 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X296 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X297 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X298 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X299 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X300 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X301 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X302 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X303 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X304 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X305 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X306 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X307 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X308 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X309 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X310 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X311 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X312 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X313 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X314 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X315 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X316 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X317 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X318 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X319 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X320 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X321 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X322 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X323 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X324 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X325 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X326 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X327 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X328 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X329 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X330 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X331 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X332 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X333 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X334 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X335 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X336 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X337 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X338 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X339 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X340 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X341 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X342 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X343 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X344 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X345 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X346 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X347 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X348 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X349 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X350 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X351 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X352 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X353 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X354 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X355 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X356 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X357 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X358 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X359 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X360 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X361 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X362 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X363 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X364 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X365 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X366 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X367 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X368 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X369 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X370 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X371 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X372 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X373 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X374 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X375 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X376 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X377 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X378 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X379 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X380 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X381 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X382 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X383 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X384 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X385 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X386 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X387 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X388 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X389 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X390 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X391 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X392 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X393 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X394 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X395 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X396 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X397 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X398 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X399 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X400 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X401 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X402 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X403 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X404 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X405 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X406 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X407 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X408 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X409 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X410 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X411 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X412 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X413 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X414 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X415 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X416 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X417 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X418 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X419 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X420 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X421 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X422 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X423 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X424 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X425 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X426 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X427 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X428 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X429 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X430 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X431 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X432 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X433 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X434 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X435 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X436 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X437 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X438 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X439 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X440 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X441 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X442 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X443 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X444 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X445 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X446 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X447 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X448 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X449 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X450 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X451 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X452 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X453 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X454 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X455 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X456 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X457 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X458 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X459 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X460 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X461 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X462 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X463 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X464 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X465 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X466 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X467 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X468 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X469 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X470 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X471 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X472 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X473 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X474 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X475 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X476 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X477 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X478 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X479 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X480 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X481 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X482 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X483 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X484 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X485 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X486 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X487 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X488 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X489 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X490 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X491 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X492 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X493 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X494 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X495 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X496 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X497 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X498 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X499 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X500 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X501 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X502 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X503 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X504 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X505 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X506 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X507 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X508 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X509 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X510 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X511 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X512 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X513 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X514 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X515 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X516 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X517 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X518 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X519 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X520 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X521 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X522 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X523 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X524 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X525 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X526 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X527 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X528 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X529 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X530 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X531 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X532 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X533 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X534 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X535 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X536 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X537 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X538 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X539 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X540 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X541 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X542 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X543 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X544 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X545 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X546 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X547 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X548 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X549 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X550 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X551 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X552 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X553 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X554 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X555 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X556 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X557 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X558 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X559 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X560 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X561 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X562 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X563 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X564 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X565 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X566 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X567 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X568 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X569 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X570 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X571 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X572 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X573 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X574 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X575 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X576 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X577 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X578 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X579 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X580 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X581 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X582 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X583 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X584 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X585 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X586 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X587 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X588 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X589 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X590 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X591 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X592 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X593 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X594 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X595 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X596 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X597 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X598 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X599 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X600 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X601 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X602 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X603 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X604 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X605 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X606 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X607 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X608 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X609 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X610 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X611 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X612 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X613 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X614 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X615 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X616 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X617 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X618 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X619 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X620 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X621 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X622 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X623 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X624 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X625 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X626 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X627 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X628 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X629 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X630 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X631 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X632 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X633 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X634 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X635 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X636 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X637 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X638 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X639 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X640 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X641 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X642 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X643 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X644 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X645 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X646 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X647 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X648 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X649 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X650 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X651 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X652 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X653 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X654 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X655 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X656 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X657 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X658 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X659 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X660 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X661 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X662 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X663 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X664 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X665 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X666 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X667 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X668 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X669 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X670 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X671 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X672 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X673 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X674 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X675 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X676 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X677 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X678 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X679 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X680 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X681 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X682 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X683 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X684 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X685 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X686 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X687 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X688 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X689 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X690 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X691 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X692 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X693 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X694 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X695 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X696 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X697 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X698 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X699 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X700 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X701 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X702 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X703 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X704 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X705 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X706 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X707 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X708 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X709 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X710 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X711 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X712 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X713 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X714 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X715 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X716 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X717 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X718 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X719 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X720 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X721 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X722 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X723 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X724 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X725 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X726 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X727 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X728 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X729 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X730 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X731 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X732 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X733 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X734 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X735 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X736 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X737 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X738 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X739 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X740 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X741 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X742 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X743 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X744 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X745 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X746 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X747 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X748 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X749 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X750 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X751 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X752 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X753 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X754 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X755 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X756 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X757 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X758 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X759 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X760 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X761 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X762 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X763 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X764 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X765 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X766 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X767 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X768 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X769 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X770 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X771 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X772 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X773 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X774 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X775 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X776 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X777 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X778 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X779 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X780 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X781 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X782 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X783 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X784 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X785 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X786 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X787 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X788 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X789 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X790 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X791 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X792 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X793 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X794 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X795 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X796 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X797 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X798 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X799 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X800 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X801 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X802 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X803 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X804 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X805 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X806 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X807 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X808 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X809 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X810 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X811 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X812 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X813 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X814 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X815 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X816 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X817 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X818 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X819 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X820 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X821 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X822 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X823 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X824 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X825 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X826 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X827 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X828 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X829 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X830 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X831 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X832 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X833 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X834 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X835 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X836 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X837 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X838 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X839 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X840 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X841 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X842 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X843 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X844 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X845 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X846 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X847 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X848 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X849 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X850 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X851 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X852 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X853 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X854 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X855 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X856 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X857 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X858 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X859 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X860 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X861 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X862 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X863 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X864 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X865 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X866 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X867 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X868 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X869 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X870 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X871 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X872 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X873 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X874 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X875 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X876 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X877 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X878 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X879 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X880 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X881 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X882 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X883 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X884 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X885 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X886 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X887 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X888 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X889 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X890 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X891 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X892 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X893 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X894 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X895 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X896 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X897 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X898 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X899 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X900 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X901 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X902 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X903 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X904 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X905 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X906 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X907 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X908 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X909 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X910 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X911 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X912 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X913 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X914 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X915 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X916 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X917 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X918 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X919 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X920 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X921 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X922 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X923 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X924 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X925 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X926 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X927 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X928 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X929 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X930 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X931 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X932 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X933 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X934 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X935 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X936 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X937 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X938 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X939 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X940 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X941 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X942 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X943 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X944 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X945 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X946 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X947 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X948 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X949 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X950 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X951 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X952 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X953 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X954 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X955 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X956 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X957 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X958 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X959 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X960 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X961 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X962 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X963 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X964 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X965 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X966 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X967 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X968 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X969 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X970 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X971 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X972 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X973 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X974 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X975 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X976 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X977 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X978 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X979 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X980 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X981 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X982 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X983 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X984 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X985 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X986 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X987 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X988 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X989 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X990 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X991 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X992 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X993 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X994 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X995 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X996 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X997 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X998 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X999 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1000 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1001 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1002 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1003 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1004 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1005 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1006 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1007 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1008 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1009 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1010 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1011 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1012 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1013 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1014 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1015 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1016 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1017 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1018 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1019 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1020 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1021 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1022 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1023 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1024 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1025 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1026 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1027 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1028 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1029 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1030 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1031 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1032 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1033 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1034 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1035 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1036 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1037 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1038 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1039 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1040 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1041 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1042 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1043 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1044 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1045 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1046 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1047 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1048 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1049 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1050 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1051 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1052 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1053 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1054 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1055 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1056 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1057 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1058 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1059 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1060 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1061 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1062 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1063 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1064 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1065 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1066 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1067 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1068 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1069 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1070 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1071 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1072 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1073 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1074 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1075 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1076 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1077 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1078 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1079 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1080 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1081 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1082 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1083 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1084 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1085 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1086 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1087 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1088 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1089 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1090 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1091 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1092 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1093 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1094 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1095 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1096 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1097 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1098 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1099 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1100 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1101 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1102 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1103 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1104 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1105 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1106 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1107 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1108 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1109 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1110 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1111 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1112 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1113 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1114 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1115 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1116 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1117 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1118 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1119 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1120 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1121 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1122 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1123 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1124 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1125 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1126 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1127 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1128 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1129 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1130 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1131 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1132 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1133 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1134 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1135 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1136 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1137 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1138 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1139 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1140 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1141 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1142 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1143 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1144 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1145 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1146 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1147 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1148 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1149 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1150 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1151 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1152 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1153 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1154 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1155 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1156 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1157 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1158 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1159 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1160 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1161 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1162 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1163 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1164 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1165 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1166 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1167 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1168 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1169 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1170 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1171 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1172 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1173 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1174 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1175 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1176 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1177 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1178 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1179 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1180 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1181 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1182 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1183 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1184 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1185 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1186 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1187 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1188 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1189 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1190 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1191 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1192 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1193 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1194 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1195 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1196 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1197 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1198 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1199 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1200 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1201 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1202 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1203 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1204 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1205 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1206 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1207 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1208 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1209 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1210 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1211 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1212 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1213 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1214 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1215 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1216 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1217 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1218 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1219 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1220 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1221 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1222 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1223 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1224 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1225 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1226 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1227 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1228 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1229 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1230 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1231 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1232 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1233 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1234 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1235 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1236 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1237 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1238 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1239 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1240 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1241 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1242 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1243 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1244 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1245 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1246 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1247 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1248 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1249 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1250 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1251 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1252 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1253 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1254 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1255 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1256 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1257 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1258 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1259 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1260 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1261 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1262 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1263 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1264 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1265 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1266 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1267 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1268 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1269 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1270 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1271 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1272 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1273 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1274 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1275 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1276 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1277 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1278 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1279 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1280 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1281 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1282 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1283 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1284 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1285 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1286 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1287 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1288 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1289 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1290 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1291 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1292 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1293 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1294 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1295 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1296 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1297 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1298 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1299 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1300 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1301 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1302 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1303 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1304 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1305 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1306 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1307 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1308 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1309 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1310 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1311 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1312 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1313 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1314 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1315 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1316 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1317 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1318 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1319 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1320 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1321 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1322 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1323 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1324 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1325 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1326 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1327 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1328 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1329 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1330 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1331 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1332 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1333 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1334 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1335 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1336 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1337 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1338 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1339 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1340 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1341 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1342 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1343 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1344 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1345 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1346 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1347 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1348 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1349 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1350 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1351 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1352 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1353 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1354 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1355 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1356 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1357 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1358 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1359 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1360 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1361 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1362 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1363 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1364 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1365 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1366 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1367 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1368 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1369 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1370 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1371 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1372 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1373 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1374 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1375 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1376 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1377 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1378 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1379 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1380 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1381 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1382 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1383 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1384 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1385 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1386 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1387 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1388 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1389 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1390 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1391 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1392 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1393 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1394 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1395 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1396 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1397 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1398 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1399 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1400 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1401 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1402 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1403 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1404 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1405 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1406 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1407 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1408 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1409 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1410 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1411 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1412 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1413 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1414 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1415 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1416 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1417 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1418 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1419 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1420 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1421 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1422 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1423 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1424 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1425 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1426 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1427 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1428 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1429 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1430 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1431 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1432 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1433 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1434 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1435 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1436 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1437 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1438 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1439 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1440 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1441 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1442 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1443 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1444 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1445 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1446 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1447 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1448 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1449 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1450 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1451 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1452 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1453 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1454 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1455 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1456 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1457 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1458 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1459 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1460 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1461 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1462 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1463 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1464 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1465 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1466 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1467 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1468 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1469 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1470 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1471 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1472 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1473 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1474 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1475 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1476 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1477 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1478 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1479 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1480 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1481 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1482 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1483 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1484 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1485 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1486 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1487 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1488 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1489 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1490 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1491 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1492 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1493 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1494 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1495 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1496 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1497 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1498 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1499 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1500 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1501 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1502 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1503 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1504 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1505 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1506 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1507 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1508 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1509 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1510 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1511 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1512 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1513 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1514 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1515 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1516 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1517 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1518 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1519 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1520 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1521 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1522 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1523 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1524 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1525 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1526 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1527 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1528 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1529 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1530 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1531 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1532 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1533 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1534 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1535 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1536 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1537 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1538 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1539 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1540 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1541 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1542 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1543 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1544 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1545 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1546 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1547 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1548 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1549 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1550 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1551 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1552 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1553 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1554 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1555 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1556 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1557 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1558 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1559 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1560 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1561 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1562 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1563 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1564 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1565 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1566 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1567 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1568 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1569 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1570 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1571 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1572 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1573 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1574 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1575 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1576 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1577 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1578 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1579 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1580 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1581 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1582 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1583 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1584 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1585 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1586 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1587 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1588 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1589 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1590 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1591 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1592 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1593 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1594 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1595 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1596 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1597 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1598 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1599 VDDIN NDRIVE VSSOUT VSSOUT sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
.ends

* expanding   symbol:  powerp.sym # of pins=3
** sym_path: /home/nikhil/Desktop/Basic_Boost_Converter/Spice_Files/powerp.sym
** sch_path: /home/nikhil/Desktop/Basic_Boost_Converter/Spice_Files/powerp.sch
.subckt powerp  Pdrive VDDIN VSSOUT
*.ipin Pdrive
*.iopin VSSOUT
*.iopin VDDIN

X0 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X2 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X3 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X4 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X5 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X6 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X7 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X8 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X9 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X10 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X11 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X12 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X13 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X14 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X15 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X16 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X17 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X18 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X19 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X20 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X21 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X22 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X23 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X24 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X25 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X26 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X27 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X28 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X29 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X30 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X31 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X32 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X33 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X34 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X35 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X36 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X37 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X38 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X39 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X40 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X41 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X42 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X43 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X44 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X45 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X46 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X47 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X48 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X49 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X50 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X51 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X52 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X53 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X54 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X55 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X56 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X57 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X58 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X59 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X60 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X61 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X62 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X63 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X64 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X65 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X66 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X67 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X68 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X69 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X70 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X71 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X72 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X73 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X74 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X75 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X76 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X77 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X78 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X79 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X80 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X81 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X82 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X83 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X84 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X85 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X86 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X87 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X88 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X89 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X90 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X91 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X92 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X93 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X94 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X95 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X96 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X97 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X98 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X99 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X100 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X101 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X102 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X103 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X104 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X105 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X106 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X107 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X108 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X109 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X110 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X111 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X112 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X113 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X114 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X115 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X116 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X117 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X118 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X119 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X120 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X121 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X122 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X123 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X124 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X125 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X126 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X127 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X128 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X129 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X130 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X131 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X132 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X133 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X134 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X135 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X136 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X137 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X138 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X139 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X140 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X141 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X142 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X143 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X144 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X145 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X146 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X147 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X148 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X149 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X150 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X151 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X152 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X153 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X154 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X155 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X156 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X157 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X158 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X159 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X160 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X161 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X162 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X163 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X164 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X165 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X166 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X167 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X168 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X169 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X170 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X171 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X172 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X173 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X174 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X175 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X176 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X177 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X178 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X179 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X180 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X181 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X182 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X183 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X184 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X185 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X186 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X187 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X188 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X189 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X190 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X191 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X192 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X193 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X194 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X195 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X196 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X197 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X198 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X199 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X200 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X201 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X202 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X203 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X204 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X205 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X206 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X207 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X208 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X209 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X210 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X211 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X212 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X213 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X214 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X215 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X216 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X217 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X218 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X219 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X220 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X221 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X222 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X223 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X224 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X225 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X226 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X227 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X228 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X229 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X230 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X231 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X232 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X233 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X234 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X235 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X236 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X237 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X238 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X239 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X240 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X241 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X242 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X243 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X244 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X245 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X246 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X247 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X248 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X249 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X250 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X251 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X252 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X253 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X254 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X255 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X256 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X257 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X258 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X259 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X260 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X261 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X262 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X263 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X264 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X265 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X266 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X267 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X268 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X269 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X270 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X271 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X272 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X273 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X274 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X275 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X276 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X277 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X278 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X279 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X280 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X281 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X282 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X283 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X284 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X285 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X286 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X287 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X288 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X289 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X290 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X291 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X292 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X293 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X294 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X295 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X296 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X297 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X298 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X299 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X300 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X301 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X302 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X303 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X304 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X305 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X306 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X307 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X308 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X309 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X310 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X311 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X312 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X313 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X314 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X315 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X316 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X317 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X318 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X319 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X320 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X321 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X322 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X323 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X324 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X325 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X326 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X327 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X328 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X329 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X330 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X331 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X332 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X333 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X334 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X335 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X336 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X337 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X338 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X339 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X340 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X341 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X342 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X343 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X344 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X345 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X346 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X347 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X348 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X349 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X350 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X351 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X352 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X353 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X354 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X355 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X356 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X357 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X358 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X359 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X360 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X361 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X362 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X363 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X364 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X365 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X366 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X367 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X368 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X369 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X370 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X371 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X372 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X373 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X374 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X375 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X376 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X377 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X378 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X379 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X380 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X381 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X382 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X383 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X384 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X385 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X386 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X387 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X388 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X389 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X390 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X391 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X392 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X393 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X394 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X395 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X396 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X397 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X398 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X399 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X400 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X401 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X402 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X403 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X404 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X405 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X406 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X407 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X408 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X409 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X410 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X411 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X412 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X413 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X414 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X415 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X416 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X417 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X418 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X419 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X420 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X421 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X422 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X423 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X424 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X425 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X426 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X427 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X428 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X429 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X430 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X431 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X432 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X433 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X434 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X435 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X436 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X437 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X438 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X439 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X440 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X441 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X442 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X443 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X444 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X445 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X446 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X447 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X448 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X449 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X450 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X451 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X452 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X453 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X454 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X455 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X456 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X457 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X458 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X459 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X460 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X461 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X462 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X463 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X464 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X465 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X466 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X467 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X468 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X469 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X470 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X471 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X472 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X473 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X474 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X475 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X476 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X477 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X478 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X479 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X480 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X481 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X482 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X483 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X484 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X485 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X486 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X487 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X488 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X489 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X490 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X491 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X492 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X493 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X494 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X495 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X496 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X497 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X498 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X499 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X500 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X501 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X502 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X503 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X504 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X505 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X506 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X507 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X508 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X509 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X510 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X511 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X512 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X513 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X514 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X515 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X516 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X517 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X518 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X519 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X520 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X521 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X522 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X523 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X524 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X525 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X526 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X527 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X528 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X529 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X530 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X531 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X532 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X533 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X534 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X535 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X536 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X537 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X538 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X539 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X540 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X541 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X542 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X543 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X544 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X545 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X546 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X547 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X548 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X549 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X550 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X551 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X552 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X553 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X554 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X555 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X556 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X557 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X558 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X559 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X560 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X561 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X562 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X563 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X564 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X565 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X566 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X567 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X568 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X569 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X570 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X571 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X572 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X573 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X574 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X575 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X576 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X577 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X578 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X579 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X580 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X581 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X582 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X583 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X584 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X585 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X586 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X587 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X588 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X589 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X590 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X591 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X592 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X593 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X594 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X595 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X596 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X597 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X598 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X599 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X600 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X601 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X602 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X603 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X604 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X605 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X606 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X607 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X608 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X609 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X610 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X611 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X612 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X613 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X614 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X615 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X616 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X617 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X618 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X619 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X620 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X621 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X622 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X623 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X624 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X625 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X626 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X627 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X628 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X629 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X630 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X631 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X632 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X633 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X634 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X635 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X636 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X637 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X638 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X639 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X640 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X641 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X642 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X643 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X644 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X645 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X646 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X647 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X648 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X649 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X650 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X651 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X652 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X653 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X654 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X655 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X656 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X657 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X658 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X659 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X660 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X661 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X662 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X663 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X664 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X665 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X666 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X667 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X668 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X669 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X670 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X671 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X672 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X673 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X674 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X675 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X676 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X677 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X678 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X679 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X680 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X681 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X682 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X683 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X684 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X685 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X686 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X687 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X688 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X689 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X690 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X691 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X692 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X693 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X694 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X695 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X696 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X697 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X698 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X699 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X700 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X701 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X702 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X703 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X704 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X705 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X706 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X707 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X708 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X709 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X710 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X711 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X712 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X713 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X714 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X715 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X716 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X717 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X718 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X719 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X720 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X721 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X722 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X723 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X724 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X725 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X726 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X727 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X728 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X729 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X730 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X731 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X732 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X733 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X734 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X735 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X736 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X737 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X738 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X739 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X740 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X741 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X742 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X743 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X744 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X745 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X746 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X747 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X748 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X749 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X750 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X751 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X752 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X753 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X754 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X755 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X756 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X757 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X758 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X759 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X760 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X761 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X762 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X763 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X764 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X765 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X766 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X767 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X768 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X769 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X770 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X771 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X772 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X773 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X774 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X775 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X776 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X777 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X778 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X779 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X780 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X781 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X782 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X783 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X784 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X785 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X786 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X787 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X788 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X789 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X790 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X791 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X792 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X793 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X794 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X795 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X796 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X797 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X798 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X799 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X800 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X801 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X802 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X803 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X804 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X805 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X806 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X807 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X808 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X809 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X810 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X811 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X812 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X813 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X814 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X815 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X816 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X817 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X818 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X819 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X820 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X821 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X822 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X823 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X824 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X825 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X826 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X827 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X828 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X829 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X830 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X831 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X832 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X833 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X834 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X835 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X836 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X837 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X838 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X839 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X840 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X841 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X842 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X843 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X844 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X845 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X846 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X847 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X848 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X849 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X850 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X851 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X852 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X853 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X854 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X855 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X856 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X857 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X858 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X859 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X860 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X861 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X862 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X863 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X864 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X865 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X866 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X867 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X868 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X869 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X870 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X871 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X872 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X873 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X874 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X875 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X876 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X877 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X878 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X879 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X880 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X881 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X882 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X883 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X884 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X885 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X886 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X887 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X888 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X889 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X890 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X891 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X892 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X893 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X894 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X895 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X896 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X897 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X898 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X899 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X900 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X901 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X902 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X903 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X904 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X905 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X906 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X907 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X908 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X909 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X910 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X911 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X912 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X913 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X914 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X915 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X916 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X917 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X918 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X919 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X920 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X921 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X922 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X923 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X924 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X925 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X926 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X927 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X928 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X929 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X930 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X931 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X932 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X933 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X934 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X935 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X936 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X937 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X938 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X939 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X940 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X941 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X942 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X943 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X944 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X945 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X946 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X947 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X948 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X949 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X950 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X951 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X952 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X953 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X954 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X955 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X956 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X957 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X958 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X959 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X960 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X961 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X962 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X963 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X964 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X965 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X966 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X967 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X968 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X969 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X970 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X971 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X972 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X973 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X974 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X975 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X976 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X977 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X978 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X979 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X980 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X981 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X982 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X983 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X984 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X985 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X986 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X987 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X988 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X989 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X990 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X991 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X992 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X993 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X994 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X995 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X996 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X997 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X998 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X999 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1000 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1001 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1002 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1003 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1004 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1005 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1006 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1007 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1008 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1009 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1010 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1011 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1012 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1013 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1014 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1015 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1016 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1017 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1018 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1019 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1020 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1021 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1022 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1023 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1024 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1025 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1026 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1027 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1028 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1029 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1030 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1031 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1032 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1033 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1034 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1035 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1036 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1037 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1038 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1039 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1040 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1041 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1042 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1043 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1044 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1045 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1046 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1047 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1048 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1049 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1050 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1051 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1052 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1053 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1054 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1055 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1056 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1057 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1058 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1059 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1060 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1061 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1062 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1063 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1064 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1065 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1066 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1067 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1068 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1069 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1070 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1071 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1072 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1073 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1074 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1075 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1076 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1077 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1078 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1079 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1080 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1081 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1082 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1083 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1084 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1085 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1086 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1087 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1088 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1089 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1090 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1091 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1092 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1093 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1094 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1095 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1096 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1097 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1098 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1099 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1100 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1101 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1102 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1103 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1104 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1105 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1106 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1107 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1108 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1109 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1110 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1111 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1112 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1113 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1114 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1115 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1116 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1117 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1118 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1119 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1120 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1121 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1122 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1123 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1124 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1125 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1126 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1127 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1128 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1129 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1130 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1131 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1132 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1133 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1134 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1135 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1136 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1137 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1138 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1139 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1140 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1141 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1142 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1143 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1144 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1145 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1146 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1147 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1148 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1149 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1150 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1151 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1152 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1153 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1154 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1155 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1156 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1157 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1158 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1159 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1160 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1161 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1162 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1163 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1164 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1165 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1166 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1167 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1168 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1169 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1170 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1171 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1172 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1173 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1174 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1175 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1176 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1177 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1178 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1179 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1180 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1181 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1182 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1183 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1184 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1185 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1186 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1187 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1188 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1189 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1190 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1191 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1192 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1193 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1194 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1195 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1196 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1197 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1198 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1199 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1200 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1201 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1202 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1203 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1204 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1205 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1206 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1207 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1208 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1209 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1210 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1211 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1212 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1213 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1214 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1215 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1216 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1217 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1218 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1219 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1220 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1221 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1222 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1223 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1224 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1225 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1226 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1227 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1228 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1229 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1230 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1231 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1232 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1233 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1234 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1235 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1236 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1237 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1238 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1239 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1240 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1241 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1242 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1243 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1244 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1245 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1246 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1247 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1248 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1249 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1250 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1251 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1252 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1253 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1254 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1255 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1256 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1257 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1258 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1259 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1260 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1261 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1262 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1263 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1264 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1265 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1266 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1267 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1268 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1269 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1270 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1271 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1272 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1273 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1274 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1275 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1276 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1277 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1278 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1279 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1280 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1281 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1282 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1283 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1284 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1285 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1286 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1287 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1288 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1289 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1290 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1291 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1292 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1293 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1294 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1295 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1296 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1297 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1298 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1299 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1300 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1301 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1302 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1303 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1304 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1305 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1306 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1307 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1308 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1309 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1310 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1311 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1312 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1313 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1314 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1315 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1316 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1317 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1318 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1319 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1320 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1321 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1322 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1323 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1324 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1325 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1326 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1327 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1328 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1329 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1330 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1331 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1332 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1333 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1334 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1335 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1336 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1337 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1338 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1339 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1340 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1341 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1342 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1343 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1344 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1345 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1346 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1347 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1348 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1349 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1350 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1351 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1352 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1353 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1354 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1355 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1356 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1357 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1358 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1359 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1360 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1361 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1362 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1363 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1364 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1365 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1366 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1367 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1368 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1369 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1370 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1371 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1372 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1373 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1374 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1375 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1376 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1377 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1378 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1379 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1380 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1381 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1382 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1383 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1384 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1385 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1386 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1387 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1388 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1389 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1390 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1391 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1392 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1393 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1394 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1395 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1396 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1397 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1398 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1399 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1400 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1401 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1402 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1403 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1404 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1405 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1406 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1407 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1408 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1409 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1410 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1411 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1412 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1413 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1414 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1415 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1416 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1417 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1418 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1419 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1420 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1421 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1422 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1423 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1424 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1425 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1426 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1427 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1428 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1429 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1430 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1431 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1432 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1433 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1434 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1435 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1436 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1437 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1438 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1439 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1440 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1441 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1442 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1443 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1444 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1445 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1446 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1447 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1448 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1449 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1450 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1451 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1452 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1453 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1454 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1455 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1456 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1457 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1458 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1459 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1460 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1461 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1462 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1463 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1464 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1465 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1466 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1467 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1468 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1469 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1470 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1471 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1472 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1473 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1474 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1475 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1476 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1477 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1478 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1479 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1480 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1481 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1482 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1483 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1484 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1485 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1486 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1487 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1488 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1489 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1490 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1491 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1492 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1493 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1494 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1495 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1496 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1497 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1498 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1499 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1500 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1501 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1502 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1503 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1504 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1505 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1506 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1507 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1508 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1509 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1510 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1511 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1512 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1513 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1514 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1515 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1516 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1517 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1518 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1519 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1520 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1521 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1522 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1523 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1524 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1525 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1526 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1527 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1528 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1529 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1530 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1531 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1532 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1533 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1534 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1535 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1536 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1537 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1538 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1539 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1540 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1541 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1542 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1543 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1544 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1545 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1546 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1547 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1548 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1549 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1550 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1551 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1552 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1553 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1554 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1555 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1556 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1557 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1558 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1559 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1560 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1561 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1562 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1563 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1564 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1565 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1566 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1567 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1568 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1569 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1570 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1571 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1572 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1573 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1574 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1575 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1576 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1577 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1578 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1579 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1580 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1581 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1582 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1583 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1584 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1585 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1586 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1587 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1588 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1589 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1590 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1591 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1592 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1593 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1594 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1595 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1596 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1597 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1598 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1599 VDDIN Pdrive VSSOUT VSSOUT sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
.ends

.GLOBAL GND
.end
