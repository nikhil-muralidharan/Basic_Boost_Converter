magic
tech sky130A
timestamp 1659421205
<< error_s >>
rect 321 280 925 359
<< nwell >>
rect -205 275 925 280
rect -205 115 405 275
<< pmoslvt >>
rect -55 145 -20 245
rect 30 145 65 245
rect 215 145 250 245
<< nmoslvt >>
rect -55 -50 -40 50
rect 90 -50 105 50
rect 235 -50 250 50
<< ndiff >>
rect -105 35 -55 50
rect -105 -35 -90 35
rect -70 -35 -55 35
rect -105 -50 -55 -35
rect -40 35 10 50
rect -40 -35 -25 35
rect -5 -35 10 35
rect -40 -50 10 -35
rect 40 35 90 50
rect 40 -35 55 35
rect 75 -35 90 35
rect 40 -50 90 -35
rect 105 35 155 50
rect 105 -35 120 35
rect 140 -35 155 35
rect 105 -50 155 -35
rect 185 35 235 50
rect 185 -35 200 35
rect 220 -35 235 35
rect 185 -50 235 -35
rect 250 35 300 50
rect 250 -35 265 35
rect 285 -35 300 35
rect 250 -50 300 -35
<< pdiff >>
rect -105 230 -55 245
rect -105 160 -90 230
rect -70 160 -55 230
rect -105 145 -55 160
rect -20 230 30 245
rect -20 160 -5 230
rect 15 160 30 230
rect -20 145 30 160
rect 65 230 115 245
rect 65 160 80 230
rect 100 160 115 230
rect 65 145 115 160
rect 165 230 215 245
rect 165 160 180 230
rect 200 160 215 230
rect 165 145 215 160
rect 250 230 300 245
rect 250 160 265 230
rect 285 160 300 230
rect 250 145 300 160
<< ndiffc >>
rect -90 -35 -70 35
rect -25 -35 -5 35
rect 55 -35 75 35
rect 120 -35 140 35
rect 200 -35 220 35
rect 265 -35 285 35
<< pdiffc >>
rect -90 160 -70 230
rect -5 160 15 230
rect 80 160 100 230
rect 180 160 200 230
rect 265 160 285 230
<< psubdiff >>
rect -185 35 -135 50
rect -185 -35 -170 35
rect -150 -35 -135 35
rect -185 -50 -135 -35
<< nsubdiff >>
rect -185 230 -135 245
rect -185 160 -170 230
rect -150 160 -135 230
rect -185 145 -135 160
<< psubdiffcont >>
rect -170 -35 -150 35
<< nsubdiffcont >>
rect -170 160 -150 230
<< poly >>
rect -55 245 -20 260
rect 30 245 65 260
rect 215 245 250 260
rect -55 130 -20 145
rect 30 130 65 145
rect 215 130 250 145
rect -55 50 -40 130
rect 50 80 65 130
rect 235 105 250 130
rect 195 95 250 105
rect 50 65 105 80
rect 195 75 205 95
rect 225 75 250 95
rect 195 65 250 75
rect 90 50 105 65
rect 235 50 250 65
rect -55 -65 -40 -50
rect 90 -65 105 -50
rect 235 -65 250 -50
rect -55 -75 -15 -65
rect -55 -95 -45 -75
rect -25 -95 -15 -75
rect -55 -105 -15 -95
rect 90 -75 130 -65
rect 90 -95 100 -75
rect 120 -95 130 -75
rect 90 -105 130 -95
<< polycont >>
rect 205 75 225 95
rect -45 -95 -25 -75
rect 100 -95 120 -75
<< locali >>
rect -180 230 -140 240
rect -180 160 -170 230
rect -150 160 -140 230
rect -180 150 -140 160
rect -100 230 -60 240
rect -100 160 -90 230
rect -70 160 -60 230
rect -100 150 -60 160
rect -15 230 25 240
rect -15 160 -5 230
rect 15 160 25 230
rect -15 150 25 160
rect 70 230 110 240
rect 70 160 80 230
rect 100 160 110 230
rect 70 150 110 160
rect 170 230 210 240
rect 170 160 180 230
rect 200 160 210 230
rect 170 150 210 160
rect 255 230 295 240
rect 255 160 265 230
rect 285 160 295 230
rect 255 150 295 160
rect 80 95 100 150
rect 195 95 235 105
rect -25 75 205 95
rect 225 75 235 95
rect -25 45 -5 75
rect 120 45 140 75
rect 195 65 235 75
rect 275 100 295 150
rect 275 80 375 100
rect 275 45 295 80
rect -180 35 -140 45
rect -180 -35 -170 35
rect -150 -35 -140 35
rect -180 -45 -140 -35
rect -100 35 -60 45
rect -100 -35 -90 35
rect -70 -35 -60 35
rect -100 -45 -60 -35
rect -35 35 5 45
rect -35 -35 -25 35
rect -5 -35 5 35
rect -35 -45 5 -35
rect 45 35 85 45
rect 45 -35 55 35
rect 75 -35 85 35
rect 45 -45 85 -35
rect 110 35 150 45
rect 110 -35 120 35
rect 140 -35 150 35
rect 110 -45 150 -35
rect 190 35 230 45
rect 190 -35 200 35
rect 220 -35 230 35
rect 190 -45 230 -35
rect 255 35 295 45
rect 255 -35 265 35
rect 285 -35 295 35
rect 255 -45 295 -35
rect 355 -65 375 80
rect -55 -75 -15 -65
rect -55 -95 -45 -75
rect -25 -95 -15 -75
rect -55 -105 -15 -95
rect 90 -75 130 -65
rect 90 -95 100 -75
rect 120 -95 130 -75
rect 355 -85 410 -65
rect 90 -105 130 -95
<< viali >>
rect -170 160 -150 230
rect -90 160 -70 230
rect 180 160 200 230
rect -170 -35 -150 35
rect -90 -35 -70 35
rect 55 -35 75 35
rect 200 -35 220 35
<< metal1 >>
rect -205 230 405 240
rect -205 160 -170 230
rect -150 160 -90 230
rect -70 160 180 230
rect 200 160 405 230
rect -205 150 405 160
rect -205 35 405 45
rect -205 -35 -170 35
rect -150 -35 -90 35
rect -70 -35 55 35
rect 75 -35 200 35
rect 220 -35 405 35
rect -205 -45 405 -35
use and_lvt  and_lvt_0
timestamp 1659421205
transform 1 0 -75 0 1 -615
box -160 0 500 405
use inverter_lvt  inverter_lvt_0
timestamp 1658301810
transform 1 0 860 0 1 -535
box -185 -80 75 300
use inverter_lvt  inverter_lvt_1
timestamp 1658301810
transform 1 0 600 0 1 -535
box -185 -80 75 300
<< labels >>
rlabel metal1 -205 195 -205 195 7 VP
port 1 w
rlabel metal1 -205 0 -205 0 7 VN
port 2 w
rlabel locali -35 -105 -35 -105 5 A
port 3 s
rlabel locali 110 -105 110 -105 5 B
port 4 s
rlabel locali 335 90 335 90 3 Y
port 5 e
<< end >>
