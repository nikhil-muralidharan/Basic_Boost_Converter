magic
tech sky130A
timestamp 1640179147
<< end >>
