magic
tech sky130A
timestamp 1658392855
<< nwell >>
rect -115 70 145 205
<< pmoslvt >>
rect 40 90 75 185
<< nmoslvt >>
rect 35 -100 50 -5
<< ndiff >>
rect -15 -20 35 -5
rect -15 -85 0 -20
rect 20 -85 35 -20
rect -15 -100 35 -85
rect 50 -20 100 -5
rect 50 -85 65 -20
rect 85 -85 100 -20
rect 50 -100 100 -85
<< pdiff >>
rect -10 170 40 185
rect -10 105 5 170
rect 25 105 40 170
rect -10 90 40 105
rect 75 170 125 185
rect 75 105 90 170
rect 110 105 125 170
rect 75 90 125 105
<< ndiffc >>
rect 0 -85 20 -20
rect 65 -85 85 -20
<< pdiffc >>
rect 5 105 25 170
rect 90 105 110 170
<< psubdiff >>
rect -95 -20 -45 -5
rect -95 -85 -80 -20
rect -60 -85 -45 -20
rect -95 -100 -45 -85
<< nsubdiff >>
rect -95 170 -45 185
rect -95 105 -80 170
rect -60 105 -45 170
rect -95 90 -45 105
<< psubdiffcont >>
rect -80 -85 -60 -20
<< nsubdiffcont >>
rect -80 105 -60 170
<< poly >>
rect 25 245 75 255
rect 25 225 35 245
rect 55 225 75 245
rect 25 216 75 225
rect 40 185 75 216
rect 40 70 75 90
rect 35 -5 50 10
rect 35 -130 50 -100
rect 10 -140 50 -130
rect 10 -160 20 -140
rect 40 -160 50 -140
rect 10 -169 50 -160
<< polycont >>
rect 35 225 55 245
rect 20 -160 40 -140
<< locali >>
rect 35 255 55 270
rect 25 245 65 255
rect 25 225 35 245
rect 55 225 65 245
rect 25 216 65 225
rect -90 170 -50 180
rect -90 105 -80 170
rect -60 105 -50 170
rect -90 95 -50 105
rect -5 170 35 180
rect -5 105 5 170
rect 25 105 35 170
rect -5 95 35 105
rect 80 170 120 180
rect 80 105 90 170
rect 110 105 120 170
rect 80 95 120 105
rect 5 35 25 95
rect 90 40 110 95
rect -115 20 25 35
rect 65 20 145 40
rect -115 15 20 20
rect 0 -10 20 15
rect 65 -10 85 20
rect -90 -20 -50 -10
rect -90 -85 -80 -20
rect -60 -85 -50 -20
rect -90 -95 -50 -85
rect -10 -20 30 -10
rect -10 -85 0 -20
rect 20 -85 30 -20
rect -10 -95 30 -85
rect 55 -20 95 -10
rect 55 -85 65 -20
rect 85 -85 95 -20
rect 55 -95 95 -85
rect 10 -140 50 -130
rect 10 -160 20 -140
rect 40 -160 50 -140
rect 10 -169 50 -160
rect 20 -185 40 -169
<< viali >>
rect -80 105 -60 170
rect 90 105 110 170
rect -80 -85 -60 -20
rect 65 -85 85 -20
<< metal1 >>
rect -115 170 145 180
rect -115 105 -80 170
rect -60 105 90 170
rect 110 105 145 170
rect -115 90 145 105
rect -115 -20 145 -10
rect -115 -85 -80 -20
rect -60 -85 65 -20
rect 85 -85 145 -20
rect -115 -95 145 -85
<< labels >>
rlabel locali 145 30 145 30 3 out
port 1 e
rlabel locali -115 25 -115 25 7 in
port 2 w
rlabel locali 45 270 45 270 1 A'
port 3 n
rlabel locali 30 -185 30 -185 5 A
port 4 s
<< end >>
