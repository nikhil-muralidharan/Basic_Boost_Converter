magic
tech sky130A
timestamp 1657124887
<< nwell >>
rect -150 85 390 280
<< pmoslvt >>
rect 0 145 35 245
rect 85 145 120 245
rect 270 145 305 245
<< nmoslvt >>
rect 0 -50 15 50
rect 145 -50 160 50
rect 290 -50 305 50
<< ndiff >>
rect -50 35 0 50
rect -50 -35 -35 35
rect -15 -35 0 35
rect -50 -50 0 -35
rect 15 35 65 50
rect 15 -35 30 35
rect 50 -35 65 35
rect 15 -50 65 -35
rect 95 35 145 50
rect 95 -35 110 35
rect 130 -35 145 35
rect 95 -50 145 -35
rect 160 35 210 50
rect 160 -35 175 35
rect 195 -35 210 35
rect 160 -50 210 -35
rect 240 35 290 50
rect 240 -35 255 35
rect 275 -35 290 35
rect 240 -50 290 -35
rect 305 35 355 50
rect 305 -35 320 35
rect 340 -35 355 35
rect 305 -50 355 -35
<< pdiff >>
rect -50 230 0 245
rect -50 160 -35 230
rect -15 160 0 230
rect -50 145 0 160
rect 35 230 85 245
rect 35 160 50 230
rect 70 160 85 230
rect 35 145 85 160
rect 120 230 170 245
rect 120 160 135 230
rect 155 160 170 230
rect 120 145 170 160
rect 220 230 270 245
rect 220 160 235 230
rect 255 160 270 230
rect 220 145 270 160
rect 305 230 355 245
rect 305 160 320 230
rect 340 160 355 230
rect 305 145 355 160
<< ndiffc >>
rect -35 -35 -15 35
rect 30 -35 50 35
rect 110 -35 130 35
rect 175 -35 195 35
rect 255 -35 275 35
rect 320 -35 340 35
<< pdiffc >>
rect -35 160 -15 230
rect 50 160 70 230
rect 135 160 155 230
rect 235 160 255 230
rect 320 160 340 230
<< psubdiff >>
rect -130 35 -80 50
rect -130 -35 -115 35
rect -95 -35 -80 35
rect -130 -50 -80 -35
<< nsubdiff >>
rect -130 230 -80 245
rect -130 160 -115 230
rect -95 160 -80 230
rect -130 145 -80 160
<< psubdiffcont >>
rect -115 -35 -95 35
<< nsubdiffcont >>
rect -115 160 -95 230
<< poly >>
rect 0 245 35 260
rect 85 245 120 260
rect 270 245 305 260
rect 0 130 35 145
rect 85 130 120 145
rect 270 130 305 145
rect 0 50 15 130
rect 105 80 120 130
rect 290 105 305 130
rect 250 95 305 105
rect 105 65 160 80
rect 250 75 260 95
rect 280 75 305 95
rect 250 65 305 75
rect 145 50 160 65
rect 290 50 305 65
rect 0 -65 15 -50
rect 145 -65 160 -50
rect 290 -65 305 -50
rect 0 -75 40 -65
rect 0 -95 10 -75
rect 30 -95 40 -75
rect 0 -105 40 -95
rect 145 -75 185 -65
rect 145 -95 155 -75
rect 175 -95 185 -75
rect 145 -105 185 -95
<< polycont >>
rect 260 75 280 95
rect 10 -95 30 -75
rect 155 -95 175 -75
<< locali >>
rect -125 230 -85 240
rect -125 160 -115 230
rect -95 160 -85 230
rect -125 150 -85 160
rect -45 230 -5 240
rect -45 160 -35 230
rect -15 160 -5 230
rect -45 150 -5 160
rect 40 230 80 240
rect 40 160 50 230
rect 70 160 80 230
rect 40 150 80 160
rect 125 230 165 240
rect 125 160 135 230
rect 155 160 165 230
rect 125 150 165 160
rect 225 230 265 240
rect 225 160 235 230
rect 255 160 265 230
rect 225 150 265 160
rect 310 230 350 240
rect 310 160 320 230
rect 340 160 350 230
rect 310 150 350 160
rect 135 95 155 150
rect 250 95 290 105
rect 30 75 260 95
rect 280 75 290 95
rect 30 45 50 75
rect 175 45 195 75
rect 250 65 290 75
rect 330 100 350 150
rect 330 80 390 100
rect 330 45 350 80
rect -125 35 -85 45
rect -125 -35 -115 35
rect -95 -35 -85 35
rect -125 -45 -85 -35
rect -45 35 -5 45
rect -45 -35 -35 35
rect -15 -35 -5 35
rect -45 -45 -5 -35
rect 20 35 60 45
rect 20 -35 30 35
rect 50 -35 60 35
rect 20 -45 60 -35
rect 100 35 140 45
rect 100 -35 110 35
rect 130 -35 140 35
rect 100 -45 140 -35
rect 165 35 205 45
rect 165 -35 175 35
rect 195 -35 205 35
rect 165 -45 205 -35
rect 245 35 285 45
rect 245 -35 255 35
rect 275 -35 285 35
rect 245 -45 285 -35
rect 310 35 350 45
rect 310 -35 320 35
rect 340 -35 350 35
rect 310 -45 350 -35
rect 0 -75 40 -65
rect 0 -95 10 -75
rect 30 -95 40 -75
rect 0 -105 40 -95
rect 145 -75 185 -65
rect 145 -95 155 -75
rect 175 -95 185 -75
rect 145 -105 185 -95
<< viali >>
rect -115 160 -95 230
rect -35 160 -15 230
rect 235 160 255 230
rect -115 -35 -95 35
rect -35 -35 -15 35
rect 110 -35 130 35
rect 255 -35 275 35
<< metal1 >>
rect -150 230 390 245
rect -150 160 -115 230
rect -95 160 -35 230
rect -15 160 235 230
rect 255 160 390 230
rect -150 145 390 160
rect -150 35 390 45
rect -150 -35 -115 35
rect -95 -35 -35 35
rect -15 -35 110 35
rect 130 -35 255 35
rect 275 -35 390 35
rect -150 -45 390 -35
<< end >>
