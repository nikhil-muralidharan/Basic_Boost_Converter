magic
tech sky130A
magscale 1 2
timestamp 1640157656
<< nmos >>
rect -15 -2000 15 2000
<< ndiff >>
rect -73 1988 -15 2000
rect -73 -1988 -61 1988
rect -27 -1988 -15 1988
rect -73 -2000 -15 -1988
rect 15 1988 73 2000
rect 15 -1988 27 1988
rect 61 -1988 73 1988
rect 15 -2000 73 -1988
<< ndiffc >>
rect -61 -1988 -27 1988
rect 27 -1988 61 1988
<< poly >>
rect -15 2000 15 2026
rect -15 -2026 15 -2000
<< locali >>
rect -61 1988 -27 2004
rect -61 -2004 -27 -1988
rect 27 1988 61 2004
rect 27 -2004 61 -1988
<< viali >>
rect -61 -1988 -27 1988
rect 27 -1988 61 1988
<< metal1 >>
rect -67 1988 -21 2000
rect -67 -1988 -61 1988
rect -27 -1988 -21 1988
rect -67 -2000 -21 -1988
rect 21 1988 67 2000
rect 21 -1988 27 1988
rect 61 -1988 67 1988
rect 21 -2000 67 -1988
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 20 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
