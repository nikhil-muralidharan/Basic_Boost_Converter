* SPICE3 file created from basic_boost_1.ext - technology: sky130A

.subckt power_nmos_2 a_1290_520# a_890_n50#
X0 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X2 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X3 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X4 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X5 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X6 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X7 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X8 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X9 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X10 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X11 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X12 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X13 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X14 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X15 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X16 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X17 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X18 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X19 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X20 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X21 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X22 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X23 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X24 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X25 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X26 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X27 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X28 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X29 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X30 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X31 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X32 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X33 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X34 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X35 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X36 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X37 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X38 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X39 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X40 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X41 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X42 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X43 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X44 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X45 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X46 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X47 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X48 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X49 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X50 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X51 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X52 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X53 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X54 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X55 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X56 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X57 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X58 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X59 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X60 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X61 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X62 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X63 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X64 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X65 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X66 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X67 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X68 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X69 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X70 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X71 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X72 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X73 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X74 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X75 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X76 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X77 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X78 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X79 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X80 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X81 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X82 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X83 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X84 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X85 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X86 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X87 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X88 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X89 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X90 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X91 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X92 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X93 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X94 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X95 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X96 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X97 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X98 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X99 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X100 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X101 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X102 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X103 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X104 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X105 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X106 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X107 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X108 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X109 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X110 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X111 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X112 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X113 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X114 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X115 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X116 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X117 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X118 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X119 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X120 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X121 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X122 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X123 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X124 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X125 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X126 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X127 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X128 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X129 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X130 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X131 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X132 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X133 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X134 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X135 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X136 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X137 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X138 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X139 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X140 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X141 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X142 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X143 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X144 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X145 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X146 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X147 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X148 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X149 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X150 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X151 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X152 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X153 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X154 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X155 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X156 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X157 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X158 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X159 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X160 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X161 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X162 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X163 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X164 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X165 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X166 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X167 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X168 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X169 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X170 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X171 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X172 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X173 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X174 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X175 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X176 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X177 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X178 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X179 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X180 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X181 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X182 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X183 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X184 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X185 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X186 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X187 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X188 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X189 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X190 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X191 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X192 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X193 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X194 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X195 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X196 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X197 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X198 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X199 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X200 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X201 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X202 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X203 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X204 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X205 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X206 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X207 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X208 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X209 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X210 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X211 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X212 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X213 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X214 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X215 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X216 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X217 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X218 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X219 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X220 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X221 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X222 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X223 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X224 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X225 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X226 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X227 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X228 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X229 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X230 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X231 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X232 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X233 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X234 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X235 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X236 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X237 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X238 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X239 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X240 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X241 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X242 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X243 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X244 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X245 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X246 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X247 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X248 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X249 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X250 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X251 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X252 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X253 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X254 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X255 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X256 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X257 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X258 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X259 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X260 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X261 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X262 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X263 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X264 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X265 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X266 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X267 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X268 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X269 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X270 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X271 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X272 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X273 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X274 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X275 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X276 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X277 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X278 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X279 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X280 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X281 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X282 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X283 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X284 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X285 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X286 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X287 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X288 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X289 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X290 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X291 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X292 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X293 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X294 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X295 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X296 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X297 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X298 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X299 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X300 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X301 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X302 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X303 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X304 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X305 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X306 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X307 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X308 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X309 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X310 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X311 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X312 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X313 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X314 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X315 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X316 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X317 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X318 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X319 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X320 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X321 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X322 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X323 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X324 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X325 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X326 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X327 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X328 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X329 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X330 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X331 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X332 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X333 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X334 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X335 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X336 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X337 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X338 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X339 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X340 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X341 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X342 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X343 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X344 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X345 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X346 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X347 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X348 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X349 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X350 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X351 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X352 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X353 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X354 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X355 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X356 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X357 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X358 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X359 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X360 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X361 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X362 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X363 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X364 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X365 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X366 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X367 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X368 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X369 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X370 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X371 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X372 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X373 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X374 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X375 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X376 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X377 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X378 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X379 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X380 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X381 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X382 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X383 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X384 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X385 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X386 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X387 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X388 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X389 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X390 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X391 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X392 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X393 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X394 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X395 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X396 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X397 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X398 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X399 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X400 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X401 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X402 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X403 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X404 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X405 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X406 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X407 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X408 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X409 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X410 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X411 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X412 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X413 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X414 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X415 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X416 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X417 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X418 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X419 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X420 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X421 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X422 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X423 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X424 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X425 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X426 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X427 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X428 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X429 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X430 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X431 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X432 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X433 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X434 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X435 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X436 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X437 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X438 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X439 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X440 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X441 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X442 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X443 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X444 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X445 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X446 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X447 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X448 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X449 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X450 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X451 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X452 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X453 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X454 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X455 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X456 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X457 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X458 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X459 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X460 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X461 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X462 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X463 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X464 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X465 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X466 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X467 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X468 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X469 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X470 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X471 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X472 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X473 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X474 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X475 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X476 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X477 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X478 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X479 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X480 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X481 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X482 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X483 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X484 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X485 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X486 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X487 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X488 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X489 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X490 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X491 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X492 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X493 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X494 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X495 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X496 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X497 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X498 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X499 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X500 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X501 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X502 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X503 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X504 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X505 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X506 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X507 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X508 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X509 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X510 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X511 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X512 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X513 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X514 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X515 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X516 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X517 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X518 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X519 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X520 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X521 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X522 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X523 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X524 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X525 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X526 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X527 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X528 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X529 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X530 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X531 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X532 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X533 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X534 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X535 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X536 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X537 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X538 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X539 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X540 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X541 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X542 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X543 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X544 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X545 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X546 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X547 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X548 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X549 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X550 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X551 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X552 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X553 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X554 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X555 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X556 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X557 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X558 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X559 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X560 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X561 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X562 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X563 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X564 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X565 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X566 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X567 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X568 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X569 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X570 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X571 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X572 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X573 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X574 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X575 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X576 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X577 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X578 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X579 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X580 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X581 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X582 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X583 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X584 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X585 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X586 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X587 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X588 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X589 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X590 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X591 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X592 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X593 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X594 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X595 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X596 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X597 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X598 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X599 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X600 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X601 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X602 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X603 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X604 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X605 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X606 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X607 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X608 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X609 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X610 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X611 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X612 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X613 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X614 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X615 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X616 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X617 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X618 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X619 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X620 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X621 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X622 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X623 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X624 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X625 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X626 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X627 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X628 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X629 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X630 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X631 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X632 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X633 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X634 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X635 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X636 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X637 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X638 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X639 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X640 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X641 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X642 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X643 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X644 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X645 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X646 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X647 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X648 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X649 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X650 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X651 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X652 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X653 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X654 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X655 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X656 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X657 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X658 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X659 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X660 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X661 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X662 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X663 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X664 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X665 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X666 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X667 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X668 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X669 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X670 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X671 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X672 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X673 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X674 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X675 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X676 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X677 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X678 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X679 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X680 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X681 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X682 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X683 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X684 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X685 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X686 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X687 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X688 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X689 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X690 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X691 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X692 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X693 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X694 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X695 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X696 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X697 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X698 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X699 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X700 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X701 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X702 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X703 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X704 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X705 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X706 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X707 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X708 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X709 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X710 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X711 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X712 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X713 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X714 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X715 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X716 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X717 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X718 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X719 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X720 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X721 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X722 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X723 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X724 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X725 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X726 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X727 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X728 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X729 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X730 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X731 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X732 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X733 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X734 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X735 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X736 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X737 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X738 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X739 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X740 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X741 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X742 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X743 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X744 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X745 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X746 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X747 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X748 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X749 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X750 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X751 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X752 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X753 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X754 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X755 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X756 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X757 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X758 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X759 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X760 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X761 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X762 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X763 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X764 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X765 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X766 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X767 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X768 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X769 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X770 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X771 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X772 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X773 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X774 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X775 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X776 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X777 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X778 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X779 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X780 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X781 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X782 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X783 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X784 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X785 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X786 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X787 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X788 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X789 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X790 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X791 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X792 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X793 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X794 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X795 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X796 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X797 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X798 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X799 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X800 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X801 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X802 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X803 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X804 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X805 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X806 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X807 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X808 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X809 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X810 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X811 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X812 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X813 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X814 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X815 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X816 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X817 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X818 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X819 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X820 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X821 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X822 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X823 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X824 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X825 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X826 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X827 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X828 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X829 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X830 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X831 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X832 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X833 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X834 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X835 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X836 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X837 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X838 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X839 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X840 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X841 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X842 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X843 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X844 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X845 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X846 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X847 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X848 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X849 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X850 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X851 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X852 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X853 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X854 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X855 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X856 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X857 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X858 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X859 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X860 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X861 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X862 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X863 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X864 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X865 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X866 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X867 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X868 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X869 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X870 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X871 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X872 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X873 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X874 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X875 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X876 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X877 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X878 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X879 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X880 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X881 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X882 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X883 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X884 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X885 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X886 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X887 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X888 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X889 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X890 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X891 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X892 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X893 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X894 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X895 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X896 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X897 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X898 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X899 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X900 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X901 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X902 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X903 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X904 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X905 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X906 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X907 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X908 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X909 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X910 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X911 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X912 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X913 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X914 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X915 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X916 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X917 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X918 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X919 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X920 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X921 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X922 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X923 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X924 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X925 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X926 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X927 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X928 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X929 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X930 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X931 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X932 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X933 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X934 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X935 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X936 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X937 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X938 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X939 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X940 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X941 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X942 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X943 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X944 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X945 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X946 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X947 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X948 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X949 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X950 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X951 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X952 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X953 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X954 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X955 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X956 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X957 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X958 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X959 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X960 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X961 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X962 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X963 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X964 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X965 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X966 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X967 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X968 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X969 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X970 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X971 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X972 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X973 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X974 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X975 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X976 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X977 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X978 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X979 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X980 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X981 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X982 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X983 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X984 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X985 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X986 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X987 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X988 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X989 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X990 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X991 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X992 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X993 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X994 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X995 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X996 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X997 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X998 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X999 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1000 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1001 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1002 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1003 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1004 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1005 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1006 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1007 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1008 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1009 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1010 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1011 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1012 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1013 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1014 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1015 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1016 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1017 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1018 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1019 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1020 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1021 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1022 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1023 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1024 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1025 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1026 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1027 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1028 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1029 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1030 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1031 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1032 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1033 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1034 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1035 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1036 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1037 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1038 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1039 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1040 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1041 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1042 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1043 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1044 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1045 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1046 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1047 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1048 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1049 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1050 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1051 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1052 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1053 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1054 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1055 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1056 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1057 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1058 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1059 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1060 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1061 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1062 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1063 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1064 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1065 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1066 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1067 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1068 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1069 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1070 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1071 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1072 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1073 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1074 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1075 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1076 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1077 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1078 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1079 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1080 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1081 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1082 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1083 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1084 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1085 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1086 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1087 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1088 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1089 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1090 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1091 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1092 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1093 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1094 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1095 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1096 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1097 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1098 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1099 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1100 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1101 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1102 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1103 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1104 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1105 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1106 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1107 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1108 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1109 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1110 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1111 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1112 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1113 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1114 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1115 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1116 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1117 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1118 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1119 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1120 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1121 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1122 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1123 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1124 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1125 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1126 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1127 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1128 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1129 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1130 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1131 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1132 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1133 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1134 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1135 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1136 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1137 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1138 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1139 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1140 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1141 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1142 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1143 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1144 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1145 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1146 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1147 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1148 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1149 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1150 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1151 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1152 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1153 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1154 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1155 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1156 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1157 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1158 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1159 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1160 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1161 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1162 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1163 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1164 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1165 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1166 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1167 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1168 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1169 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1170 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1171 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1172 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1173 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1174 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1175 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1176 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1177 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1178 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1179 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1180 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1181 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1182 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1183 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1184 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1185 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1186 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1187 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1188 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1189 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1190 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1191 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1192 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1193 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1194 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1195 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1196 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1197 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1198 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1199 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1200 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1201 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1202 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1203 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1204 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1205 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1206 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1207 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1208 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1209 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1210 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1211 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1212 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1213 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1214 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1215 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1216 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1217 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1218 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1219 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1220 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1221 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1222 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1223 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1224 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1225 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1226 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1227 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1228 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1229 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1230 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1231 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1232 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1233 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1234 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1235 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1236 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1237 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1238 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1239 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1240 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1241 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1242 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1243 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1244 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1245 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1246 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1247 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1248 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1249 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1250 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1251 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1252 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1253 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1254 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1255 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1256 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1257 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1258 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1259 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1260 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1261 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1262 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1263 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1264 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1265 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1266 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1267 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1268 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1269 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1270 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1271 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1272 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1273 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1274 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1275 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1276 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1277 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1278 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1279 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1280 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1281 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1282 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1283 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1284 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1285 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1286 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1287 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1288 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1289 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1290 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1291 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1292 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1293 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1294 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1295 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1296 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1297 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1298 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1299 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1300 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1301 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1302 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1303 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1304 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1305 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1306 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1307 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1308 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1309 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1310 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1311 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1312 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1313 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1314 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1315 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1316 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1317 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1318 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1319 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1320 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1321 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1322 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1323 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1324 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1325 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1326 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1327 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1328 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1329 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1330 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1331 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1332 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1333 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1334 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1335 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1336 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1337 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1338 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1339 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1340 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1341 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1342 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1343 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1344 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1345 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1346 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1347 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1348 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1349 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1350 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1351 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1352 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1353 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1354 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1355 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1356 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1357 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1358 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1359 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1360 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1361 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1362 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1363 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1364 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1365 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1366 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1367 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1368 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1369 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1370 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1371 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1372 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1373 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1374 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1375 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1376 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1377 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1378 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1379 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1380 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1381 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1382 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1383 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1384 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1385 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1386 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1387 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1388 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1389 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1390 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1391 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1392 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1393 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1394 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1395 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1396 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1397 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1398 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1399 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1400 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1401 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1402 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1403 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1404 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1405 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1406 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1407 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1408 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1409 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1410 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1411 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1412 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1413 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1414 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1415 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1416 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1417 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1418 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1419 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1420 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1421 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1422 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1423 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1424 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1425 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1426 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1427 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1428 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1429 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1430 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1431 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1432 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1433 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1434 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1435 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1436 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1437 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1438 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1439 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1440 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1441 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1442 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1443 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1444 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1445 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1446 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1447 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1448 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1449 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1450 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1451 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1452 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1453 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1454 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1455 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1456 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1457 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1458 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1459 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1460 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1461 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1462 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1463 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1464 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1465 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1466 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1467 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1468 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1469 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1470 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1471 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1472 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1473 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1474 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1475 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1476 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1477 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1478 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1479 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1480 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1481 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1482 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1483 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1484 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1485 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1486 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1487 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1488 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1489 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1490 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1491 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1492 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1493 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1494 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1495 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1496 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1497 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1498 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1499 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1500 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1501 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1502 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1503 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1504 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1505 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1506 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1507 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1508 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1509 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1510 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1511 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1512 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1513 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1514 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1515 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1516 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1517 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1518 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1519 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1520 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1521 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1522 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1523 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1524 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1525 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1526 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1527 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1528 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1529 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1530 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1531 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1532 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1533 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1534 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1535 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1536 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1537 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1538 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1539 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1540 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1541 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1542 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1543 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1544 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1545 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1546 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1547 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1548 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1549 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1550 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1551 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1552 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1553 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1554 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1555 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1556 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1557 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1558 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1559 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1560 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1561 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1562 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1563 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1564 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1565 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1566 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1567 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1568 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1569 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1570 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1571 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1572 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1573 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1574 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1575 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1576 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1577 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1578 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1579 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1580 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1581 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1582 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1583 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1584 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1585 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1586 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1587 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1588 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1589 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1590 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1591 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1592 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1593 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1594 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1595 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1596 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1597 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1598 a_1290_520# a_1490_400# a_1520_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1599 a_1520_520# a_1490_400# a_1290_520# a_890_n50# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
C0 a_1290_520# a_1520_520# 5592.90fF
C1 a_1490_400# a_1290_520# 34.67fF
C2 a_1490_400# a_1520_520# 34.67fF
C3 a_1520_520# a_890_n50# 596.95fF
C4 a_1290_520# a_890_n50# 667.21fF
C5 a_1490_400# a_890_n50# 955.88fF
.ends

.subckt power_pmos_2 a_1290_520# VSUBS w_n690_n690#
X0 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=1.6848e+16p pd=3.536e+10u as=1.6848e+16p ps=3.536e+10u w=2.025e+07u l=150000u
X1 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X2 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X3 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X4 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X5 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X6 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X7 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X8 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X9 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X10 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X11 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X12 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X13 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X14 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X15 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X16 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X17 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X18 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X19 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X20 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X21 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X22 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X23 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X24 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X25 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X26 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X27 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X28 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X29 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X30 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X31 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X32 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X33 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X34 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X35 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X36 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X37 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X38 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X39 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X40 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X41 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X42 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X43 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X44 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X45 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X46 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X47 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X48 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X49 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X50 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X51 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X52 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X53 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X54 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X55 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X56 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X57 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X58 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X59 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X60 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X61 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X62 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X63 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X64 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X65 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X66 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X67 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X68 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X69 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X70 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X71 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X72 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X73 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X74 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X75 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X76 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X77 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X78 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X79 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X80 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X81 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X82 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X83 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X84 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X85 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X86 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X87 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X88 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X89 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X90 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X91 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X92 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X93 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X94 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X95 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X96 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X97 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X98 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X99 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X100 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X101 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X102 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X103 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X104 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X105 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X106 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X107 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X108 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X109 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X110 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X111 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X112 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X113 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X114 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X115 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X116 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X117 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X118 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X119 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X120 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X121 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X122 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X123 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X124 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X125 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X126 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X127 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X128 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X129 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X130 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X131 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X132 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X133 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X134 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X135 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X136 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X137 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X138 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X139 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X140 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X141 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X142 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X143 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X144 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X145 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X146 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X147 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X148 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X149 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X150 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X151 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X152 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X153 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X154 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X155 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X156 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X157 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X158 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X159 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X160 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X161 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X162 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X163 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X164 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X165 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X166 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X167 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X168 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X169 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X170 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X171 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X172 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X173 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X174 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X175 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X176 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X177 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X178 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X179 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X180 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X181 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X182 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X183 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X184 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X185 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X186 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X187 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X188 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X189 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X190 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X191 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X192 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X193 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X194 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X195 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X196 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X197 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X198 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X199 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X200 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X201 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X202 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X203 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X204 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X205 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X206 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X207 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X208 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X209 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X210 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X211 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X212 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X213 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X214 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X215 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X216 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X217 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X218 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X219 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X220 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X221 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X222 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X223 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X224 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X225 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X226 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X227 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X228 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X229 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X230 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X231 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X232 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X233 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X234 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X235 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X236 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X237 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X238 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X239 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X240 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X241 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X242 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X243 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X244 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X245 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X246 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X247 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X248 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X249 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X250 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X251 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X252 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X253 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X254 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X255 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X256 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X257 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X258 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X259 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X260 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X261 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X262 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X263 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X264 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X265 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X266 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X267 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X268 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X269 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X270 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X271 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X272 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X273 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X274 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X275 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X276 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X277 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X278 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X279 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X280 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X281 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X282 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X283 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X284 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X285 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X286 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X287 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X288 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X289 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X290 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X291 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X292 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X293 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X294 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X295 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X296 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X297 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X298 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X299 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X300 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X301 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X302 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X303 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X304 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X305 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X306 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X307 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X308 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X309 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X310 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X311 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X312 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X313 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X314 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X315 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X316 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X317 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X318 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X319 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X320 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X321 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X322 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X323 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X324 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X325 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X326 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X327 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X328 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X329 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X330 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X331 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X332 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X333 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X334 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X335 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X336 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X337 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X338 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X339 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X340 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X341 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X342 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X343 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X344 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X345 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X346 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X347 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X348 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X349 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X350 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X351 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X352 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X353 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X354 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X355 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X356 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X357 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X358 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X359 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X360 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X361 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X362 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X363 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X364 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X365 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X366 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X367 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X368 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X369 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X370 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X371 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X372 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X373 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X374 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X375 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X376 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X377 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X378 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X379 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X380 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X381 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X382 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X383 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X384 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X385 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X386 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X387 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X388 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X389 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X390 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X391 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X392 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X393 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X394 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X395 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X396 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X397 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X398 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X399 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X400 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X401 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X402 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X403 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X404 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X405 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X406 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X407 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X408 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X409 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X410 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X411 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X412 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X413 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X414 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X415 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X416 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X417 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X418 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X419 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X420 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X421 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X422 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X423 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X424 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X425 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X426 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X427 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X428 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X429 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X430 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X431 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X432 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X433 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X434 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X435 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X436 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X437 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X438 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X439 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X440 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X441 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X442 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X443 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X444 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X445 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X446 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X447 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X448 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X449 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X450 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X451 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X452 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X453 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X454 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X455 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X456 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X457 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X458 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X459 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X460 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X461 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X462 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X463 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X464 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X465 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X466 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X467 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X468 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X469 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X470 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X471 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X472 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X473 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X474 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X475 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X476 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X477 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X478 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X479 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X480 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X481 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X482 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X483 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X484 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X485 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X486 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X487 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X488 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X489 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X490 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X491 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X492 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X493 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X494 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X495 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X496 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X497 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X498 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X499 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X500 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X501 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X502 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X503 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X504 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X505 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X506 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X507 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X508 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X509 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X510 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X511 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X512 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X513 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X514 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X515 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X516 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X517 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X518 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X519 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X520 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X521 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X522 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X523 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X524 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X525 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X526 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X527 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X528 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X529 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X530 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X531 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X532 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X533 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X534 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X535 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X536 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X537 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X538 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X539 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X540 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X541 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X542 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X543 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X544 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X545 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X546 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X547 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X548 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X549 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X550 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X551 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X552 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X553 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X554 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X555 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X556 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X557 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X558 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X559 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X560 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X561 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X562 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X563 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X564 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X565 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X566 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X567 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X568 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X569 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X570 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X571 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X572 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X573 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X574 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X575 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X576 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X577 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X578 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X579 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X580 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X581 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X582 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X583 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X584 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X585 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X586 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X587 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X588 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X589 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X590 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X591 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X592 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X593 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X594 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X595 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X596 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X597 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X598 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X599 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X600 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X601 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X602 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X603 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X604 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X605 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X606 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X607 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X608 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X609 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X610 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X611 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X612 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X613 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X614 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X615 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X616 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X617 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X618 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X619 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X620 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X621 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X622 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X623 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X624 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X625 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X626 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X627 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X628 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X629 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X630 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X631 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X632 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X633 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X634 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X635 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X636 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X637 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X638 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X639 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X640 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X641 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X642 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X643 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X644 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X645 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X646 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X647 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X648 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X649 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X650 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X651 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X652 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X653 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X654 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X655 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X656 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X657 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X658 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X659 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X660 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X661 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X662 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X663 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X664 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X665 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X666 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X667 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X668 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X669 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X670 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X671 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X672 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X673 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X674 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X675 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X676 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X677 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X678 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X679 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X680 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X681 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X682 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X683 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X684 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X685 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X686 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X687 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X688 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X689 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X690 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X691 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X692 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X693 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X694 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X695 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X696 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X697 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X698 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X699 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X700 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X701 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X702 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X703 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X704 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X705 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X706 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X707 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X708 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X709 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X710 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X711 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X712 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X713 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X714 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X715 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X716 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X717 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X718 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X719 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X720 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X721 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X722 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X723 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X724 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X725 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X726 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X727 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X728 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X729 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X730 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X731 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X732 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X733 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X734 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X735 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X736 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X737 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X738 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X739 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X740 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X741 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X742 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X743 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X744 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X745 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X746 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X747 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X748 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X749 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X750 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X751 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X752 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X753 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X754 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X755 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X756 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X757 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X758 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X759 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X760 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X761 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X762 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X763 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X764 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X765 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X766 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X767 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X768 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X769 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X770 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X771 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X772 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X773 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X774 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X775 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X776 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X777 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X778 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X779 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X780 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X781 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X782 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X783 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X784 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X785 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X786 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X787 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X788 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X789 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X790 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X791 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X792 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X793 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X794 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X795 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X796 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X797 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X798 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X799 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X800 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X801 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X802 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X803 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X804 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X805 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X806 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X807 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X808 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X809 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X810 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X811 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X812 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X813 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X814 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X815 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X816 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X817 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X818 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X819 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X820 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X821 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X822 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X823 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X824 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X825 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X826 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X827 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X828 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X829 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X830 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X831 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X832 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X833 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X834 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X835 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X836 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X837 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X838 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X839 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X840 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X841 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X842 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X843 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X844 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X845 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X846 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X847 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X848 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X849 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X850 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X851 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X852 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X853 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X854 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X855 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X856 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X857 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X858 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X859 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X860 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X861 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X862 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X863 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X864 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X865 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X866 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X867 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X868 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X869 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X870 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X871 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X872 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X873 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X874 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X875 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X876 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X877 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X878 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X879 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X880 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X881 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X882 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X883 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X884 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X885 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X886 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X887 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X888 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X889 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X890 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X891 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X892 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X893 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X894 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X895 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X896 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X897 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X898 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X899 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X900 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X901 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X902 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X903 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X904 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X905 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X906 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X907 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X908 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X909 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X910 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X911 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X912 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X913 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X914 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X915 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X916 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X917 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X918 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X919 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X920 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X921 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X922 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X923 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X924 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X925 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X926 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X927 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X928 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X929 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X930 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X931 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X932 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X933 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X934 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X935 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X936 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X937 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X938 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X939 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X940 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X941 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X942 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X943 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X944 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X945 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X946 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X947 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X948 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X949 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X950 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X951 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X952 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X953 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X954 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X955 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X956 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X957 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X958 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X959 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X960 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X961 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X962 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X963 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X964 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X965 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X966 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X967 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X968 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X969 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X970 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X971 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X972 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X973 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X974 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X975 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X976 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X977 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X978 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X979 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X980 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X981 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X982 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X983 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X984 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X985 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X986 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X987 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X988 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X989 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X990 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X991 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X992 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X993 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X994 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X995 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X996 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X997 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X998 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X999 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1000 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1001 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1002 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1003 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1004 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1005 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1006 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1007 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1008 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1009 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1010 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1011 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1012 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1013 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1014 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1015 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1016 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1017 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1018 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1019 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1020 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1021 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1022 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1023 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1024 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1025 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1026 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1027 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1028 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1029 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1030 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1031 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1032 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1033 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1034 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1035 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1036 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1037 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1038 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1039 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1040 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1041 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1042 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1043 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1044 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1045 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1046 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1047 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1048 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1049 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1050 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1051 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1052 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1053 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1054 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1055 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1056 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1057 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1058 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1059 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1060 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1061 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1062 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1063 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1064 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1065 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1066 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1067 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1068 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1069 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1070 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1071 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1072 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1073 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1074 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1075 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1076 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1077 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1078 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1079 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1080 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1081 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1082 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1083 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1084 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1085 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1086 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1087 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1088 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1089 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1090 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1091 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1092 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1093 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1094 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1095 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1096 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1097 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1098 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1099 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1100 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1101 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1102 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1103 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1104 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1105 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1106 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1107 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1108 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1109 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1110 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1111 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1112 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1113 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1114 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1115 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1116 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1117 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1118 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1119 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1120 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1121 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1122 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1123 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1124 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1125 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1126 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1127 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1128 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1129 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1130 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1131 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1132 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1133 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1134 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1135 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1136 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1137 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1138 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1139 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1140 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1141 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1142 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1143 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1144 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1145 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1146 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1147 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1148 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1149 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1150 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1151 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1152 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1153 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1154 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1155 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1156 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1157 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1158 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1159 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1160 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1161 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1162 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1163 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1164 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1165 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1166 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1167 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1168 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1169 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1170 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1171 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1172 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1173 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1174 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1175 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1176 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1177 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1178 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1179 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1180 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1181 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1182 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1183 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1184 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1185 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1186 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1187 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1188 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1189 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1190 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1191 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1192 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1193 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1194 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1195 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1196 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1197 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1198 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1199 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1200 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1201 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1202 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1203 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1204 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1205 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1206 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1207 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1208 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1209 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1210 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1211 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1212 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1213 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1214 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1215 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1216 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1217 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1218 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1219 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1220 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1221 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1222 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1223 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1224 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1225 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1226 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1227 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1228 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1229 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1230 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1231 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1232 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1233 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1234 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1235 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1236 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1237 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1238 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1239 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1240 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1241 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1242 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1243 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1244 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1245 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1246 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1247 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1248 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1249 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1250 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1251 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1252 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1253 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1254 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1255 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1256 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1257 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1258 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1259 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1260 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1261 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1262 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1263 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1264 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1265 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1266 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1267 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1268 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1269 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1270 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1271 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1272 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1273 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1274 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1275 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1276 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1277 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1278 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1279 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1280 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1281 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1282 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1283 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1284 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1285 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1286 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1287 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1288 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1289 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1290 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1291 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1292 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1293 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1294 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1295 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1296 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1297 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1298 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1299 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1300 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1301 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1302 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1303 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1304 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1305 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1306 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1307 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1308 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1309 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1310 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1311 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1312 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1313 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1314 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1315 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1316 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1317 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1318 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1319 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1320 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1321 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1322 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1323 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1324 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1325 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1326 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1327 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1328 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1329 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1330 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1331 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1332 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1333 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1334 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1335 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1336 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1337 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1338 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1339 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1340 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1341 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1342 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1343 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1344 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1345 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1346 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1347 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1348 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1349 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1350 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1351 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1352 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1353 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1354 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1355 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1356 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1357 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1358 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1359 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1360 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1361 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1362 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1363 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1364 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1365 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1366 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1367 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1368 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1369 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1370 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1371 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1372 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1373 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1374 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1375 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1376 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1377 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1378 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1379 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1380 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1381 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1382 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1383 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1384 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1385 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1386 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1387 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1388 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1389 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1390 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1391 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1392 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1393 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1394 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1395 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1396 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1397 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1398 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1399 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1400 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1401 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1402 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1403 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1404 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1405 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1406 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1407 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1408 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1409 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1410 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1411 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1412 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1413 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1414 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1415 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1416 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1417 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1418 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1419 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1420 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1421 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1422 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1423 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1424 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1425 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1426 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1427 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1428 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1429 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1430 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1431 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1432 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1433 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1434 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1435 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1436 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1437 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1438 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1439 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1440 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1441 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1442 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1443 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1444 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1445 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1446 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1447 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1448 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1449 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1450 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1451 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1452 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1453 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1454 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1455 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1456 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1457 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1458 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1459 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1460 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1461 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1462 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1463 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1464 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1465 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1466 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1467 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1468 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1469 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1470 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1471 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1472 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1473 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1474 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1475 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1476 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1477 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1478 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1479 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1480 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1481 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1482 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1483 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1484 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1485 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1486 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1487 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1488 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1489 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1490 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1491 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1492 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1493 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1494 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1495 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1496 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1497 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1498 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1499 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1500 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1501 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1502 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1503 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1504 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1505 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1506 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1507 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1508 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1509 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1510 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1511 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1512 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1513 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1514 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1515 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1516 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1517 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1518 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1519 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1520 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1521 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1522 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1523 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1524 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1525 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1526 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1527 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1528 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1529 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1530 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1531 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1532 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1533 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1534 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1535 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1536 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1537 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1538 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1539 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1540 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1541 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1542 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1543 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1544 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1545 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1546 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1547 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1548 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1549 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1550 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1551 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1552 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1553 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1554 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1555 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1556 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1557 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1558 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1559 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1560 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1561 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1562 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1563 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1564 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1565 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1566 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1567 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1568 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1569 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1570 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1571 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1572 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1573 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1574 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1575 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1576 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1577 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1578 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1579 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1580 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1581 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1582 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1583 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1584 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1585 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1586 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1587 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1588 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1589 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1590 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1591 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1592 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1593 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1594 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1595 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1596 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1597 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1598 a_1290_520# a_1490_400# a_1520_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
X1599 a_1520_520# a_1490_400# a_1290_520# w_n690_n690# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.025e+07u l=150000u
C0 a_1490_400# a_1290_520# 34.67fF
C1 a_1290_520# a_1520_520# 5592.75fF
C2 a_1490_400# a_1520_520# 34.67fF
C3 a_1520_520# w_n690_n690# 594.77fF
C4 a_1290_520# w_n690_n690# 663.53fF
C5 a_1490_400# w_n690_n690# 955.97fF
.ends

.subckt basic_boost_1 Drain_inductor
Xpower_nmos_2_0 Drain_inductor VSUBS power_nmos_2
Xpower_pmos_2_0 Drain_inductor VSUBS w_n690_n690# power_pmos_2
C0 power_pmos_2_0/a_1520_520# power_pmos_2_0/w_n690_n690# 281.33fF **FLOATING
C1 power_pmos_2_0/a_1490_400# power_pmos_2_0/w_n690_n690# 871.06fF **FLOATING
C2 power_nmos_2_0/a_1520_520# power_pmos_2_0/w_n690_n690# 596.95fF **FLOATING
C3 Drain_inductor power_pmos_2_0/w_n690_n690# 951.76fF
C4 power_nmos_2_0/a_1490_400# power_pmos_2_0/w_n690_n690# 955.88fF **FLOATING
.ends

