magic
tech sky130A
timestamp 1659699307
<< nwell >>
rect -545 955 -535 990
rect -565 865 -535 955
rect -545 830 -535 865
rect -1475 460 0 510
rect -1475 440 -390 460
rect -1475 325 -450 440
rect -385 325 0 460
rect -1475 285 0 325
<< pmoslvt >>
rect -580 340 -545 440
<< nmoslvt >>
rect -460 665 -445 765
<< ndiff >>
rect -510 750 -460 765
rect -510 680 -495 750
rect -475 680 -460 750
rect -510 665 -460 680
rect -445 750 -395 765
rect -445 680 -430 750
rect -410 680 -395 750
rect -445 665 -395 680
<< pdiff >>
rect -630 425 -580 440
rect -630 355 -615 425
rect -595 355 -580 425
rect -630 340 -580 355
rect -545 425 -495 440
rect -545 355 -530 425
rect -510 355 -495 425
rect -545 340 -495 355
<< ndiffc >>
rect -495 680 -475 750
rect -430 680 -410 750
<< pdiffc >>
rect -615 355 -595 425
rect -530 355 -510 425
<< poly >>
rect -460 810 -420 820
rect -460 790 -450 810
rect -430 790 -420 810
rect -460 780 -420 790
rect -460 765 -445 780
rect -460 650 -445 665
rect -1320 485 -1280 495
rect -1320 465 -1310 485
rect -1290 465 -1280 485
rect -1320 455 -1280 465
rect -585 485 -545 495
rect -585 465 -575 485
rect -555 465 -545 485
rect -585 455 -545 465
rect -580 440 -545 455
rect -580 325 -545 340
<< polycont >>
rect -450 790 -430 810
rect -1310 465 -1290 485
rect -575 465 -555 485
<< xpolycontact >>
rect -1360 1040 -1325 1260
rect -1360 630 -1325 850
rect -1195 1040 -1160 1260
rect -1195 630 -1160 850
<< xpolyres >>
rect -1360 850 -1325 1040
rect -1195 850 -1160 1040
<< locali >>
rect -1325 1040 -1195 1260
rect -1475 630 -1360 850
rect -1275 590 -1250 1040
rect -460 810 -420 820
rect -460 790 -450 810
rect -430 790 -420 810
rect -460 780 -420 790
rect -1160 670 -1040 760
rect -505 750 -465 760
rect -505 680 -495 750
rect -475 680 -465 750
rect -505 670 -465 680
rect -440 750 -400 760
rect -440 680 -430 750
rect -410 680 -400 750
rect -440 670 -400 680
rect -1075 610 -895 650
rect -560 625 -540 650
rect -430 625 -410 670
rect -1075 590 -1040 610
rect -560 605 -410 625
rect -1275 560 -1040 590
rect -460 575 -440 605
rect -470 535 -430 575
rect -1320 485 -1280 495
rect -1320 465 -1310 485
rect -1290 465 -1280 485
rect -1320 455 -1280 465
rect -585 485 -545 495
rect -585 465 -575 485
rect -555 465 -545 485
rect -585 455 -545 465
rect -625 425 -585 435
rect -625 355 -615 425
rect -595 355 -585 425
rect -625 345 -585 355
rect -540 425 -500 435
rect -540 355 -530 425
rect -510 355 -500 425
rect -540 345 -500 355
rect -530 295 -510 345
rect -655 275 -510 295
rect -460 190 -440 535
rect -1215 110 -1065 130
rect -655 40 -635 110
rect -655 20 -470 40
rect -75 -25 -55 0
rect 250 -25 270 10
rect -75 -45 270 -25
<< viali >>
rect -495 680 -475 750
rect -615 355 -595 425
<< metal1 >>
rect -565 865 -535 955
rect -585 670 -550 760
rect -545 750 -335 760
rect -545 680 -495 750
rect -475 680 -335 750
rect -545 670 -335 680
rect -630 425 -470 435
rect -630 355 -615 425
rect -595 355 -470 425
rect -630 345 -470 355
rect -625 150 -605 190
rect -670 60 -470 150
use comparator_lvt_otg  comparator_lvt_otg_0
timestamp 1659595967
transform 1 0 140 0 1 335
box -140 -335 470 175
use inverter_lvt_otg  inverter_lvt_otg_0
timestamp 1658301810
transform 1 0 -1290 0 1 170
box -185 -80 75 300
use inverter_lvt_otg  inverter_lvt_otg_1
timestamp 1658301810
transform 1 0 -620 0 1 690
box -185 -80 75 300
use inverter_lvt_otg  inverter_lvt_otg_2
timestamp 1658301810
transform 1 0 -880 0 1 690
box -185 -80 75 300
use or_lvt_otg  or_lvt_otg_0
timestamp 1659683504
transform 1 0 -1010 0 1 195
box -205 -105 405 280
use trgate_lvt_otg  trgate_lvt_otg_0
timestamp 1659695591
transform 1 0 -95 0 1 175
box -375 -175 95 320
<< labels >>
rlabel space -1475 120 -1475 120 7 Pdriveb
rlabel space -900 90 -900 90 5 ZCD
rlabel locali -440 820 -440 820 1 C1
<< end >>
