magic
tech sky130A
timestamp 1660760131
<< nwell >>
rect -535 345 2690 415
rect -535 220 125 345
rect 385 220 2690 345
<< pmoslvt >>
rect -380 250 -345 350
rect -180 250 -145 350
<< nmoslvt >>
rect -380 5 -365 105
rect -315 5 -300 105
rect -65 5 -50 105
rect 0 5 15 105
rect -315 -220 -300 -120
rect -65 -220 -50 -120
<< ndiff >>
rect -430 90 -380 105
rect -430 20 -415 90
rect -395 20 -380 90
rect -430 5 -380 20
rect -365 90 -315 105
rect -365 20 -350 90
rect -330 20 -315 90
rect -365 5 -315 20
rect -300 90 -250 105
rect -300 20 -285 90
rect -265 20 -250 90
rect -300 5 -250 20
rect -115 90 -65 105
rect -115 20 -100 90
rect -80 20 -65 90
rect -115 5 -65 20
rect -50 90 0 105
rect -50 20 -35 90
rect -15 20 0 90
rect -50 5 0 20
rect 15 90 65 105
rect 15 20 30 90
rect 50 20 65 90
rect 15 5 65 20
rect -365 -135 -315 -120
rect -365 -205 -350 -135
rect -330 -205 -315 -135
rect -365 -220 -315 -205
rect -300 -135 -250 -120
rect -300 -205 -285 -135
rect -265 -205 -250 -135
rect -300 -220 -250 -205
rect -115 -135 -65 -120
rect -115 -205 -100 -135
rect -80 -205 -65 -135
rect -115 -220 -65 -205
rect -50 -135 0 -120
rect -50 -205 -35 -135
rect -15 -205 0 -135
rect -50 -220 0 -205
<< pdiff >>
rect -430 335 -380 350
rect -430 265 -415 335
rect -395 265 -380 335
rect -430 250 -380 265
rect -345 335 -295 350
rect -345 265 -330 335
rect -310 265 -295 335
rect -345 250 -295 265
rect -230 335 -180 350
rect -230 265 -215 335
rect -195 265 -180 335
rect -230 250 -180 265
rect -145 335 -95 350
rect -145 265 -130 335
rect -110 265 -95 335
rect -145 250 -95 265
<< ndiffc >>
rect -415 20 -395 90
rect -350 20 -330 90
rect -285 20 -265 90
rect -100 20 -80 90
rect -35 20 -15 90
rect 30 20 50 90
rect -350 -205 -330 -135
rect -285 -205 -265 -135
rect -100 -205 -80 -135
rect -35 -205 -15 -135
<< pdiffc >>
rect -415 265 -395 335
rect -330 265 -310 335
rect -215 265 -195 335
rect -130 265 -110 335
<< psubdiff >>
rect -515 -135 -465 -120
rect -515 -205 -500 -135
rect -480 -205 -465 -135
rect -515 -220 -465 -205
<< nsubdiff >>
rect -515 335 -465 350
rect -515 265 -500 335
rect -480 265 -465 335
rect -515 250 -465 265
<< psubdiffcont >>
rect -500 -205 -480 -135
<< nsubdiffcont >>
rect -500 265 -480 335
<< poly >>
rect -380 395 -340 405
rect -380 375 -370 395
rect -350 375 -340 395
rect -380 365 -340 375
rect -185 395 -145 405
rect -185 375 -175 395
rect -155 375 -145 395
rect -185 365 -145 375
rect -380 350 -345 365
rect -180 350 -145 365
rect -380 235 -345 250
rect -180 235 -145 250
rect -380 105 -365 125
rect -315 105 -300 125
rect -65 105 -50 125
rect 0 105 15 125
rect -380 -10 -365 5
rect -410 -20 -365 -10
rect -410 -40 -400 -20
rect -380 -40 -365 -20
rect -410 -50 -365 -40
rect -315 -10 -300 5
rect -65 -10 -50 5
rect -315 -20 -270 -10
rect -315 -40 -300 -20
rect -280 -40 -270 -20
rect -315 -50 -270 -40
rect -95 -20 -50 -10
rect -95 -40 -85 -20
rect -65 -40 -50 -20
rect -95 -50 -50 -40
rect 0 -10 15 5
rect 0 -20 45 -10
rect 0 -40 15 -20
rect 35 -40 45 -20
rect 0 -50 45 -40
rect -315 -120 -300 -100
rect -65 -120 -50 -100
rect -315 -235 -300 -220
rect -65 -235 -50 -220
rect -340 -245 -300 -235
rect -340 -265 -330 -245
rect -310 -265 -300 -245
rect -340 -275 -300 -265
rect -90 -245 -50 -235
rect -90 -265 -80 -245
rect -60 -265 -50 -245
rect -90 -275 -50 -265
<< polycont >>
rect -370 375 -350 395
rect -175 375 -155 395
rect -400 -40 -380 -20
rect -300 -40 -280 -20
rect -85 -40 -65 -20
rect 15 -40 35 -20
rect -330 -265 -310 -245
rect -80 -265 -60 -245
<< locali >>
rect -380 395 -145 405
rect -380 375 -370 395
rect -350 375 -175 395
rect -155 375 -145 395
rect -380 365 -145 375
rect -330 345 -310 365
rect -510 335 -470 345
rect -510 265 -500 335
rect -480 265 -470 335
rect -510 255 -470 265
rect -425 335 -385 345
rect -425 265 -415 335
rect -395 265 -385 335
rect -425 255 -385 265
rect -340 335 -300 345
rect -340 265 -330 335
rect -310 265 -300 335
rect -340 255 -300 265
rect -225 335 -185 345
rect -225 265 -215 335
rect -195 265 -185 335
rect -225 255 -185 265
rect -140 335 -100 345
rect -140 265 -130 335
rect -110 265 -100 335
rect -140 255 -100 265
rect -330 220 -310 255
rect -130 220 -110 255
rect -415 200 -310 220
rect -285 200 50 220
rect -415 180 -375 200
rect -415 160 -405 180
rect -385 160 -375 180
rect -415 150 -375 160
rect -415 100 -395 150
rect -285 100 -265 200
rect -120 165 -80 175
rect -120 145 -110 165
rect -90 145 -80 165
rect -120 135 -80 145
rect -100 100 -80 135
rect 30 100 50 200
rect -425 90 -385 100
rect -425 20 -415 90
rect -395 20 -385 90
rect -425 10 -385 20
rect -360 90 -320 100
rect -360 20 -350 90
rect -330 20 -320 90
rect -360 10 -320 20
rect -295 90 -255 100
rect -295 20 -285 90
rect -265 20 -255 90
rect -295 10 -255 20
rect -110 90 -70 100
rect -110 20 -100 90
rect -80 20 -70 90
rect -110 10 -70 20
rect -45 90 -5 100
rect -45 20 -35 90
rect -15 20 -5 90
rect -45 10 -5 20
rect 20 90 60 100
rect 20 20 30 90
rect 50 20 60 90
rect 20 10 60 20
rect 1540 65 1580 135
rect 1540 45 1550 65
rect 1570 45 1580 65
rect -410 -20 -370 -10
rect -410 -40 -400 -20
rect -380 -40 -370 -20
rect -410 -50 -370 -40
rect -400 -70 -380 -50
rect -425 -90 -380 -70
rect -510 -135 -470 -125
rect -510 -205 -500 -135
rect -480 -205 -470 -135
rect -510 -215 -470 -205
rect -425 -270 -405 -90
rect -350 -125 -330 10
rect -310 -20 -270 -10
rect -95 -20 -55 -10
rect -310 -40 -300 -20
rect -280 -40 -270 -20
rect -310 -50 -270 -40
rect -160 -40 -85 -20
rect -65 -40 -55 -20
rect -300 -70 -280 -50
rect -300 -90 -215 -70
rect -360 -135 -320 -125
rect -360 -205 -350 -135
rect -330 -205 -320 -135
rect -360 -215 -320 -205
rect -295 -135 -255 -125
rect -295 -205 -285 -135
rect -265 -205 -255 -135
rect -295 -215 -255 -205
rect -340 -245 -300 -235
rect -340 -265 -330 -245
rect -310 -265 -300 -245
rect -340 -275 -300 -265
rect -235 -275 -215 -90
rect -160 -275 -140 -40
rect -95 -50 -55 -40
rect -35 -125 -15 10
rect 5 -20 45 -10
rect 5 -40 15 -20
rect 35 -40 45 -20
rect 5 -50 45 -40
rect 15 -70 35 -50
rect 1540 -60 1580 45
rect 15 -90 75 -70
rect -110 -135 -70 -125
rect -110 -205 -100 -135
rect -80 -205 -70 -135
rect -110 -215 -70 -205
rect -45 -135 -5 -125
rect -45 -205 -35 -135
rect -15 -205 -5 -135
rect -45 -215 -5 -205
rect -90 -245 -50 -235
rect -90 -265 -80 -245
rect -60 -265 -50 -245
rect -90 -275 -50 -265
rect 55 -275 75 -90
rect 645 -255 795 -235
rect 1260 -255 1465 -235
rect 1920 -255 2010 -235
<< viali >>
rect -500 265 -480 335
rect -415 265 -395 335
rect -215 265 -195 335
rect -405 160 -385 180
rect -110 145 -90 165
rect 30 20 50 90
rect 1550 45 1570 65
rect -500 -205 -480 -135
rect -285 -205 -265 -135
<< metal1 >>
rect -535 335 125 345
rect -535 265 -500 335
rect -480 265 -415 335
rect -395 265 -215 335
rect -195 265 125 335
rect -535 255 125 265
rect 1255 255 1260 345
rect 1910 255 1940 345
rect -415 180 -80 190
rect -415 160 -405 180
rect -385 165 -80 180
rect -385 160 -110 165
rect -415 150 -110 160
rect -120 145 -110 150
rect -90 145 -80 165
rect -120 135 -80 145
rect -425 10 -250 100
rect -115 90 1580 100
rect -115 20 30 90
rect 50 65 1580 90
rect 50 45 1550 65
rect 1570 45 1580 65
rect 50 20 1580 45
rect -115 10 1580 20
rect -535 -135 125 -125
rect -535 -205 -500 -135
rect -480 -205 -285 -135
rect -265 -205 125 -135
rect -535 -215 125 -205
rect 1250 -215 1270 -125
rect 1890 -215 1935 -125
use and_lvt_mroat  and_lvt_mroat_0
timestamp 1660758955
transform 1 0 1420 0 1 0
box -160 -275 500 405
use inverter_lvt_mroat  inverter_lvt_mroat_0
timestamp 1660757217
transform 1 0 310 0 1 80
box -185 -355 75 300
use inverter_lvt_mroat  inverter_lvt_mroat_1
timestamp 1660757217
transform 1 0 570 0 1 80
box -185 -355 75 300
use or_lvt_mroat  or_lvt_mroat_0
timestamp 1660758149
transform 1 0 850 0 1 105
box -205 -380 410 280
use sr_latch_lvt_mroat  sr_latch_lvt_mroat_0
timestamp 1660760052
transform -1 0 2420 0 1 130
box -280 -405 505 240
<< labels >>
rlabel metal1 -535 305 -535 305 7 VP
rlabel metal1 -535 -175 -535 -175 7 VN
rlabel locali -415 -270 -415 -270 5 Vref
rlabel locali -320 -275 -320 -275 5 Vbias1
rlabel locali -225 -275 -225 -275 5 Vsen
rlabel locali -150 -275 -150 -275 5 Vsen_DC
rlabel locali -70 -275 -70 -275 1 Vbias2
rlabel space -95 -285 -95 -285 5 Vofb
rlabel space 275 -275 275 -275 5 Pdriveb
rlabel space 960 -275 960 -275 5 ZCD
rlabel space 2200 -275 2200 -275 5 CLK
<< end >>
