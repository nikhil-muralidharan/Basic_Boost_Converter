magic
tech sky130A
timestamp 1641716213
<< nwell >>
rect -1065 10070 3300 12545
rect -1070 9900 3300 10070
<< pmos >>
rect -320 10245 -305 12270
rect -205 10245 -190 12270
rect -90 10245 -75 12270
rect 25 10245 40 12270
rect 140 10245 155 12270
rect 255 10245 270 12270
rect 370 10245 385 12270
rect 485 10245 500 12270
rect 600 10245 615 12270
rect 715 10245 730 12270
rect 830 10245 845 12270
rect 945 10245 960 12270
rect 1060 10245 1075 12270
rect 1175 10245 1190 12270
rect 1290 10245 1305 12270
rect 1405 10245 1420 12270
rect 1520 10245 1535 12270
rect 1635 10245 1650 12270
rect 1750 10245 1765 12270
rect 1865 10245 1880 12270
rect 1980 10245 1995 12270
rect 2095 10245 2110 12270
rect 2210 10245 2225 12270
rect 2325 10245 2340 12270
rect 2440 10245 2455 12270
<< pdiff >>
rect -420 12235 -320 12270
rect -420 12195 -390 12235
rect -350 12195 -320 12235
rect -420 12155 -320 12195
rect -420 12115 -390 12155
rect -350 12115 -320 12155
rect -420 12075 -320 12115
rect -420 12035 -390 12075
rect -350 12035 -320 12075
rect -420 11995 -320 12035
rect -420 11955 -390 11995
rect -350 11955 -320 11995
rect -420 11915 -320 11955
rect -420 11875 -390 11915
rect -350 11875 -320 11915
rect -420 11835 -320 11875
rect -420 11795 -390 11835
rect -350 11795 -320 11835
rect -420 11755 -320 11795
rect -420 11715 -390 11755
rect -350 11715 -320 11755
rect -420 11675 -320 11715
rect -420 11635 -390 11675
rect -350 11635 -320 11675
rect -420 11595 -320 11635
rect -420 11555 -390 11595
rect -350 11555 -320 11595
rect -420 11515 -320 11555
rect -420 11475 -390 11515
rect -350 11475 -320 11515
rect -420 11435 -320 11475
rect -420 11395 -390 11435
rect -350 11395 -320 11435
rect -420 11355 -320 11395
rect -420 11315 -390 11355
rect -350 11315 -320 11355
rect -420 11275 -320 11315
rect -420 11235 -390 11275
rect -350 11235 -320 11275
rect -420 11195 -320 11235
rect -420 11155 -390 11195
rect -350 11155 -320 11195
rect -420 11115 -320 11155
rect -420 11075 -390 11115
rect -350 11075 -320 11115
rect -420 11035 -320 11075
rect -420 10995 -390 11035
rect -350 10995 -320 11035
rect -420 10955 -320 10995
rect -420 10915 -390 10955
rect -350 10915 -320 10955
rect -420 10875 -320 10915
rect -420 10835 -390 10875
rect -350 10835 -320 10875
rect -420 10795 -320 10835
rect -420 10755 -390 10795
rect -350 10755 -320 10795
rect -420 10715 -320 10755
rect -420 10675 -390 10715
rect -350 10675 -320 10715
rect -420 10635 -320 10675
rect -420 10595 -390 10635
rect -350 10595 -320 10635
rect -420 10555 -320 10595
rect -420 10515 -390 10555
rect -350 10515 -320 10555
rect -420 10475 -320 10515
rect -420 10435 -390 10475
rect -350 10435 -320 10475
rect -420 10395 -320 10435
rect -420 10355 -390 10395
rect -350 10355 -320 10395
rect -420 10315 -320 10355
rect -420 10275 -390 10315
rect -350 10275 -320 10315
rect -420 10245 -320 10275
rect -305 12235 -205 12270
rect -305 12195 -275 12235
rect -235 12195 -205 12235
rect -305 12155 -205 12195
rect -305 12115 -275 12155
rect -235 12115 -205 12155
rect -305 12075 -205 12115
rect -305 12035 -275 12075
rect -235 12035 -205 12075
rect -305 11995 -205 12035
rect -305 11955 -275 11995
rect -235 11955 -205 11995
rect -305 11915 -205 11955
rect -305 11875 -275 11915
rect -235 11875 -205 11915
rect -305 11835 -205 11875
rect -305 11795 -275 11835
rect -235 11795 -205 11835
rect -305 11755 -205 11795
rect -305 11715 -275 11755
rect -235 11715 -205 11755
rect -305 11675 -205 11715
rect -305 11635 -275 11675
rect -235 11635 -205 11675
rect -305 11595 -205 11635
rect -305 11555 -275 11595
rect -235 11555 -205 11595
rect -305 11515 -205 11555
rect -305 11475 -275 11515
rect -235 11475 -205 11515
rect -305 11435 -205 11475
rect -305 11395 -275 11435
rect -235 11395 -205 11435
rect -305 11355 -205 11395
rect -305 11315 -275 11355
rect -235 11315 -205 11355
rect -305 11275 -205 11315
rect -305 11235 -275 11275
rect -235 11235 -205 11275
rect -305 11195 -205 11235
rect -305 11155 -275 11195
rect -235 11155 -205 11195
rect -305 11115 -205 11155
rect -305 11075 -275 11115
rect -235 11075 -205 11115
rect -305 11035 -205 11075
rect -305 10995 -275 11035
rect -235 10995 -205 11035
rect -305 10955 -205 10995
rect -305 10915 -275 10955
rect -235 10915 -205 10955
rect -305 10875 -205 10915
rect -305 10835 -275 10875
rect -235 10835 -205 10875
rect -305 10795 -205 10835
rect -305 10755 -275 10795
rect -235 10755 -205 10795
rect -305 10715 -205 10755
rect -305 10675 -275 10715
rect -235 10675 -205 10715
rect -305 10635 -205 10675
rect -305 10595 -275 10635
rect -235 10595 -205 10635
rect -305 10555 -205 10595
rect -305 10515 -275 10555
rect -235 10515 -205 10555
rect -305 10475 -205 10515
rect -305 10435 -275 10475
rect -235 10435 -205 10475
rect -305 10395 -205 10435
rect -305 10355 -275 10395
rect -235 10355 -205 10395
rect -305 10315 -205 10355
rect -305 10275 -275 10315
rect -235 10275 -205 10315
rect -305 10245 -205 10275
rect -190 12235 -90 12270
rect -190 12195 -160 12235
rect -120 12195 -90 12235
rect -190 12155 -90 12195
rect -190 12115 -160 12155
rect -120 12115 -90 12155
rect -190 12075 -90 12115
rect -190 12035 -160 12075
rect -120 12035 -90 12075
rect -190 11995 -90 12035
rect -190 11955 -160 11995
rect -120 11955 -90 11995
rect -190 11915 -90 11955
rect -190 11875 -160 11915
rect -120 11875 -90 11915
rect -190 11835 -90 11875
rect -190 11795 -160 11835
rect -120 11795 -90 11835
rect -190 11755 -90 11795
rect -190 11715 -160 11755
rect -120 11715 -90 11755
rect -190 11675 -90 11715
rect -190 11635 -160 11675
rect -120 11635 -90 11675
rect -190 11595 -90 11635
rect -190 11555 -160 11595
rect -120 11555 -90 11595
rect -190 11515 -90 11555
rect -190 11475 -160 11515
rect -120 11475 -90 11515
rect -190 11435 -90 11475
rect -190 11395 -160 11435
rect -120 11395 -90 11435
rect -190 11355 -90 11395
rect -190 11315 -160 11355
rect -120 11315 -90 11355
rect -190 11275 -90 11315
rect -190 11235 -160 11275
rect -120 11235 -90 11275
rect -190 11195 -90 11235
rect -190 11155 -160 11195
rect -120 11155 -90 11195
rect -190 11115 -90 11155
rect -190 11075 -160 11115
rect -120 11075 -90 11115
rect -190 11035 -90 11075
rect -190 10995 -160 11035
rect -120 10995 -90 11035
rect -190 10955 -90 10995
rect -190 10915 -160 10955
rect -120 10915 -90 10955
rect -190 10875 -90 10915
rect -190 10835 -160 10875
rect -120 10835 -90 10875
rect -190 10795 -90 10835
rect -190 10755 -160 10795
rect -120 10755 -90 10795
rect -190 10715 -90 10755
rect -190 10675 -160 10715
rect -120 10675 -90 10715
rect -190 10635 -90 10675
rect -190 10595 -160 10635
rect -120 10595 -90 10635
rect -190 10555 -90 10595
rect -190 10515 -160 10555
rect -120 10515 -90 10555
rect -190 10475 -90 10515
rect -190 10435 -160 10475
rect -120 10435 -90 10475
rect -190 10395 -90 10435
rect -190 10355 -160 10395
rect -120 10355 -90 10395
rect -190 10315 -90 10355
rect -190 10275 -160 10315
rect -120 10275 -90 10315
rect -190 10245 -90 10275
rect -75 12235 25 12270
rect -75 12195 -45 12235
rect -5 12195 25 12235
rect -75 12155 25 12195
rect -75 12115 -45 12155
rect -5 12115 25 12155
rect -75 12075 25 12115
rect -75 12035 -45 12075
rect -5 12035 25 12075
rect -75 11995 25 12035
rect -75 11955 -45 11995
rect -5 11955 25 11995
rect -75 11915 25 11955
rect -75 11875 -45 11915
rect -5 11875 25 11915
rect -75 11835 25 11875
rect -75 11795 -45 11835
rect -5 11795 25 11835
rect -75 11755 25 11795
rect -75 11715 -45 11755
rect -5 11715 25 11755
rect -75 11675 25 11715
rect -75 11635 -45 11675
rect -5 11635 25 11675
rect -75 11595 25 11635
rect -75 11555 -45 11595
rect -5 11555 25 11595
rect -75 11515 25 11555
rect -75 11475 -45 11515
rect -5 11475 25 11515
rect -75 11435 25 11475
rect -75 11395 -45 11435
rect -5 11395 25 11435
rect -75 11355 25 11395
rect -75 11315 -45 11355
rect -5 11315 25 11355
rect -75 11275 25 11315
rect -75 11235 -45 11275
rect -5 11235 25 11275
rect -75 11195 25 11235
rect -75 11155 -45 11195
rect -5 11155 25 11195
rect -75 11115 25 11155
rect -75 11075 -45 11115
rect -5 11075 25 11115
rect -75 11035 25 11075
rect -75 10995 -45 11035
rect -5 10995 25 11035
rect -75 10955 25 10995
rect -75 10915 -45 10955
rect -5 10915 25 10955
rect -75 10875 25 10915
rect -75 10835 -45 10875
rect -5 10835 25 10875
rect -75 10795 25 10835
rect -75 10755 -45 10795
rect -5 10755 25 10795
rect -75 10715 25 10755
rect -75 10675 -45 10715
rect -5 10675 25 10715
rect -75 10635 25 10675
rect -75 10595 -45 10635
rect -5 10595 25 10635
rect -75 10555 25 10595
rect -75 10515 -45 10555
rect -5 10515 25 10555
rect -75 10475 25 10515
rect -75 10435 -45 10475
rect -5 10435 25 10475
rect -75 10395 25 10435
rect -75 10355 -45 10395
rect -5 10355 25 10395
rect -75 10315 25 10355
rect -75 10275 -45 10315
rect -5 10275 25 10315
rect -75 10245 25 10275
rect 40 12235 140 12270
rect 40 12195 70 12235
rect 110 12195 140 12235
rect 40 12155 140 12195
rect 40 12115 70 12155
rect 110 12115 140 12155
rect 40 12075 140 12115
rect 40 12035 70 12075
rect 110 12035 140 12075
rect 40 11995 140 12035
rect 40 11955 70 11995
rect 110 11955 140 11995
rect 40 11915 140 11955
rect 40 11875 70 11915
rect 110 11875 140 11915
rect 40 11835 140 11875
rect 40 11795 70 11835
rect 110 11795 140 11835
rect 40 11755 140 11795
rect 40 11715 70 11755
rect 110 11715 140 11755
rect 40 11675 140 11715
rect 40 11635 70 11675
rect 110 11635 140 11675
rect 40 11595 140 11635
rect 40 11555 70 11595
rect 110 11555 140 11595
rect 40 11515 140 11555
rect 40 11475 70 11515
rect 110 11475 140 11515
rect 40 11435 140 11475
rect 40 11395 70 11435
rect 110 11395 140 11435
rect 40 11355 140 11395
rect 40 11315 70 11355
rect 110 11315 140 11355
rect 40 11275 140 11315
rect 40 11235 70 11275
rect 110 11235 140 11275
rect 40 11195 140 11235
rect 40 11155 70 11195
rect 110 11155 140 11195
rect 40 11115 140 11155
rect 40 11075 70 11115
rect 110 11075 140 11115
rect 40 11035 140 11075
rect 40 10995 70 11035
rect 110 10995 140 11035
rect 40 10955 140 10995
rect 40 10915 70 10955
rect 110 10915 140 10955
rect 40 10875 140 10915
rect 40 10835 70 10875
rect 110 10835 140 10875
rect 40 10795 140 10835
rect 40 10755 70 10795
rect 110 10755 140 10795
rect 40 10715 140 10755
rect 40 10675 70 10715
rect 110 10675 140 10715
rect 40 10635 140 10675
rect 40 10595 70 10635
rect 110 10595 140 10635
rect 40 10555 140 10595
rect 40 10515 70 10555
rect 110 10515 140 10555
rect 40 10475 140 10515
rect 40 10435 70 10475
rect 110 10435 140 10475
rect 40 10395 140 10435
rect 40 10355 70 10395
rect 110 10355 140 10395
rect 40 10315 140 10355
rect 40 10275 70 10315
rect 110 10275 140 10315
rect 40 10245 140 10275
rect 155 12235 255 12270
rect 155 12195 185 12235
rect 225 12195 255 12235
rect 155 12155 255 12195
rect 155 12115 185 12155
rect 225 12115 255 12155
rect 155 12075 255 12115
rect 155 12035 185 12075
rect 225 12035 255 12075
rect 155 11995 255 12035
rect 155 11955 185 11995
rect 225 11955 255 11995
rect 155 11915 255 11955
rect 155 11875 185 11915
rect 225 11875 255 11915
rect 155 11835 255 11875
rect 155 11795 185 11835
rect 225 11795 255 11835
rect 155 11755 255 11795
rect 155 11715 185 11755
rect 225 11715 255 11755
rect 155 11675 255 11715
rect 155 11635 185 11675
rect 225 11635 255 11675
rect 155 11595 255 11635
rect 155 11555 185 11595
rect 225 11555 255 11595
rect 155 11515 255 11555
rect 155 11475 185 11515
rect 225 11475 255 11515
rect 155 11435 255 11475
rect 155 11395 185 11435
rect 225 11395 255 11435
rect 155 11355 255 11395
rect 155 11315 185 11355
rect 225 11315 255 11355
rect 155 11275 255 11315
rect 155 11235 185 11275
rect 225 11235 255 11275
rect 155 11195 255 11235
rect 155 11155 185 11195
rect 225 11155 255 11195
rect 155 11115 255 11155
rect 155 11075 185 11115
rect 225 11075 255 11115
rect 155 11035 255 11075
rect 155 10995 185 11035
rect 225 10995 255 11035
rect 155 10955 255 10995
rect 155 10915 185 10955
rect 225 10915 255 10955
rect 155 10875 255 10915
rect 155 10835 185 10875
rect 225 10835 255 10875
rect 155 10795 255 10835
rect 155 10755 185 10795
rect 225 10755 255 10795
rect 155 10715 255 10755
rect 155 10675 185 10715
rect 225 10675 255 10715
rect 155 10635 255 10675
rect 155 10595 185 10635
rect 225 10595 255 10635
rect 155 10555 255 10595
rect 155 10515 185 10555
rect 225 10515 255 10555
rect 155 10475 255 10515
rect 155 10435 185 10475
rect 225 10435 255 10475
rect 155 10395 255 10435
rect 155 10355 185 10395
rect 225 10355 255 10395
rect 155 10315 255 10355
rect 155 10275 185 10315
rect 225 10275 255 10315
rect 155 10245 255 10275
rect 270 12235 370 12270
rect 270 12195 300 12235
rect 340 12195 370 12235
rect 270 12155 370 12195
rect 270 12115 300 12155
rect 340 12115 370 12155
rect 270 12075 370 12115
rect 270 12035 300 12075
rect 340 12035 370 12075
rect 270 11995 370 12035
rect 270 11955 300 11995
rect 340 11955 370 11995
rect 270 11915 370 11955
rect 270 11875 300 11915
rect 340 11875 370 11915
rect 270 11835 370 11875
rect 270 11795 300 11835
rect 340 11795 370 11835
rect 270 11755 370 11795
rect 270 11715 300 11755
rect 340 11715 370 11755
rect 270 11675 370 11715
rect 270 11635 300 11675
rect 340 11635 370 11675
rect 270 11595 370 11635
rect 270 11555 300 11595
rect 340 11555 370 11595
rect 270 11515 370 11555
rect 270 11475 300 11515
rect 340 11475 370 11515
rect 270 11435 370 11475
rect 270 11395 300 11435
rect 340 11395 370 11435
rect 270 11355 370 11395
rect 270 11315 300 11355
rect 340 11315 370 11355
rect 270 11275 370 11315
rect 270 11235 300 11275
rect 340 11235 370 11275
rect 270 11195 370 11235
rect 270 11155 300 11195
rect 340 11155 370 11195
rect 270 11115 370 11155
rect 270 11075 300 11115
rect 340 11075 370 11115
rect 270 11035 370 11075
rect 270 10995 300 11035
rect 340 10995 370 11035
rect 270 10955 370 10995
rect 270 10915 300 10955
rect 340 10915 370 10955
rect 270 10875 370 10915
rect 270 10835 300 10875
rect 340 10835 370 10875
rect 270 10795 370 10835
rect 270 10755 300 10795
rect 340 10755 370 10795
rect 270 10715 370 10755
rect 270 10675 300 10715
rect 340 10675 370 10715
rect 270 10635 370 10675
rect 270 10595 300 10635
rect 340 10595 370 10635
rect 270 10555 370 10595
rect 270 10515 300 10555
rect 340 10515 370 10555
rect 270 10475 370 10515
rect 270 10435 300 10475
rect 340 10435 370 10475
rect 270 10395 370 10435
rect 270 10355 300 10395
rect 340 10355 370 10395
rect 270 10315 370 10355
rect 270 10275 300 10315
rect 340 10275 370 10315
rect 270 10245 370 10275
rect 385 12235 485 12270
rect 385 12195 415 12235
rect 455 12195 485 12235
rect 385 12155 485 12195
rect 385 12115 415 12155
rect 455 12115 485 12155
rect 385 12075 485 12115
rect 385 12035 415 12075
rect 455 12035 485 12075
rect 385 11995 485 12035
rect 385 11955 415 11995
rect 455 11955 485 11995
rect 385 11915 485 11955
rect 385 11875 415 11915
rect 455 11875 485 11915
rect 385 11835 485 11875
rect 385 11795 415 11835
rect 455 11795 485 11835
rect 385 11755 485 11795
rect 385 11715 415 11755
rect 455 11715 485 11755
rect 385 11675 485 11715
rect 385 11635 415 11675
rect 455 11635 485 11675
rect 385 11595 485 11635
rect 385 11555 415 11595
rect 455 11555 485 11595
rect 385 11515 485 11555
rect 385 11475 415 11515
rect 455 11475 485 11515
rect 385 11435 485 11475
rect 385 11395 415 11435
rect 455 11395 485 11435
rect 385 11355 485 11395
rect 385 11315 415 11355
rect 455 11315 485 11355
rect 385 11275 485 11315
rect 385 11235 415 11275
rect 455 11235 485 11275
rect 385 11195 485 11235
rect 385 11155 415 11195
rect 455 11155 485 11195
rect 385 11115 485 11155
rect 385 11075 415 11115
rect 455 11075 485 11115
rect 385 11035 485 11075
rect 385 10995 415 11035
rect 455 10995 485 11035
rect 385 10955 485 10995
rect 385 10915 415 10955
rect 455 10915 485 10955
rect 385 10875 485 10915
rect 385 10835 415 10875
rect 455 10835 485 10875
rect 385 10795 485 10835
rect 385 10755 415 10795
rect 455 10755 485 10795
rect 385 10715 485 10755
rect 385 10675 415 10715
rect 455 10675 485 10715
rect 385 10635 485 10675
rect 385 10595 415 10635
rect 455 10595 485 10635
rect 385 10555 485 10595
rect 385 10515 415 10555
rect 455 10515 485 10555
rect 385 10475 485 10515
rect 385 10435 415 10475
rect 455 10435 485 10475
rect 385 10395 485 10435
rect 385 10355 415 10395
rect 455 10355 485 10395
rect 385 10315 485 10355
rect 385 10275 415 10315
rect 455 10275 485 10315
rect 385 10245 485 10275
rect 500 12235 600 12270
rect 500 12195 530 12235
rect 570 12195 600 12235
rect 500 12155 600 12195
rect 500 12115 530 12155
rect 570 12115 600 12155
rect 500 12075 600 12115
rect 500 12035 530 12075
rect 570 12035 600 12075
rect 500 11995 600 12035
rect 500 11955 530 11995
rect 570 11955 600 11995
rect 500 11915 600 11955
rect 500 11875 530 11915
rect 570 11875 600 11915
rect 500 11835 600 11875
rect 500 11795 530 11835
rect 570 11795 600 11835
rect 500 11755 600 11795
rect 500 11715 530 11755
rect 570 11715 600 11755
rect 500 11675 600 11715
rect 500 11635 530 11675
rect 570 11635 600 11675
rect 500 11595 600 11635
rect 500 11555 530 11595
rect 570 11555 600 11595
rect 500 11515 600 11555
rect 500 11475 530 11515
rect 570 11475 600 11515
rect 500 11435 600 11475
rect 500 11395 530 11435
rect 570 11395 600 11435
rect 500 11355 600 11395
rect 500 11315 530 11355
rect 570 11315 600 11355
rect 500 11275 600 11315
rect 500 11235 530 11275
rect 570 11235 600 11275
rect 500 11195 600 11235
rect 500 11155 530 11195
rect 570 11155 600 11195
rect 500 11115 600 11155
rect 500 11075 530 11115
rect 570 11075 600 11115
rect 500 11035 600 11075
rect 500 10995 530 11035
rect 570 10995 600 11035
rect 500 10955 600 10995
rect 500 10915 530 10955
rect 570 10915 600 10955
rect 500 10875 600 10915
rect 500 10835 530 10875
rect 570 10835 600 10875
rect 500 10795 600 10835
rect 500 10755 530 10795
rect 570 10755 600 10795
rect 500 10715 600 10755
rect 500 10675 530 10715
rect 570 10675 600 10715
rect 500 10635 600 10675
rect 500 10595 530 10635
rect 570 10595 600 10635
rect 500 10555 600 10595
rect 500 10515 530 10555
rect 570 10515 600 10555
rect 500 10475 600 10515
rect 500 10435 530 10475
rect 570 10435 600 10475
rect 500 10395 600 10435
rect 500 10355 530 10395
rect 570 10355 600 10395
rect 500 10315 600 10355
rect 500 10275 530 10315
rect 570 10275 600 10315
rect 500 10245 600 10275
rect 615 12235 715 12270
rect 615 12195 645 12235
rect 685 12195 715 12235
rect 615 12155 715 12195
rect 615 12115 645 12155
rect 685 12115 715 12155
rect 615 12075 715 12115
rect 615 12035 645 12075
rect 685 12035 715 12075
rect 615 11995 715 12035
rect 615 11955 645 11995
rect 685 11955 715 11995
rect 615 11915 715 11955
rect 615 11875 645 11915
rect 685 11875 715 11915
rect 615 11835 715 11875
rect 615 11795 645 11835
rect 685 11795 715 11835
rect 615 11755 715 11795
rect 615 11715 645 11755
rect 685 11715 715 11755
rect 615 11675 715 11715
rect 615 11635 645 11675
rect 685 11635 715 11675
rect 615 11595 715 11635
rect 615 11555 645 11595
rect 685 11555 715 11595
rect 615 11515 715 11555
rect 615 11475 645 11515
rect 685 11475 715 11515
rect 615 11435 715 11475
rect 615 11395 645 11435
rect 685 11395 715 11435
rect 615 11355 715 11395
rect 615 11315 645 11355
rect 685 11315 715 11355
rect 615 11275 715 11315
rect 615 11235 645 11275
rect 685 11235 715 11275
rect 615 11195 715 11235
rect 615 11155 645 11195
rect 685 11155 715 11195
rect 615 11115 715 11155
rect 615 11075 645 11115
rect 685 11075 715 11115
rect 615 11035 715 11075
rect 615 10995 645 11035
rect 685 10995 715 11035
rect 615 10955 715 10995
rect 615 10915 645 10955
rect 685 10915 715 10955
rect 615 10875 715 10915
rect 615 10835 645 10875
rect 685 10835 715 10875
rect 615 10795 715 10835
rect 615 10755 645 10795
rect 685 10755 715 10795
rect 615 10715 715 10755
rect 615 10675 645 10715
rect 685 10675 715 10715
rect 615 10635 715 10675
rect 615 10595 645 10635
rect 685 10595 715 10635
rect 615 10555 715 10595
rect 615 10515 645 10555
rect 685 10515 715 10555
rect 615 10475 715 10515
rect 615 10435 645 10475
rect 685 10435 715 10475
rect 615 10395 715 10435
rect 615 10355 645 10395
rect 685 10355 715 10395
rect 615 10315 715 10355
rect 615 10275 645 10315
rect 685 10275 715 10315
rect 615 10245 715 10275
rect 730 12235 830 12270
rect 730 12195 760 12235
rect 800 12195 830 12235
rect 730 12155 830 12195
rect 730 12115 760 12155
rect 800 12115 830 12155
rect 730 12075 830 12115
rect 730 12035 760 12075
rect 800 12035 830 12075
rect 730 11995 830 12035
rect 730 11955 760 11995
rect 800 11955 830 11995
rect 730 11915 830 11955
rect 730 11875 760 11915
rect 800 11875 830 11915
rect 730 11835 830 11875
rect 730 11795 760 11835
rect 800 11795 830 11835
rect 730 11755 830 11795
rect 730 11715 760 11755
rect 800 11715 830 11755
rect 730 11675 830 11715
rect 730 11635 760 11675
rect 800 11635 830 11675
rect 730 11595 830 11635
rect 730 11555 760 11595
rect 800 11555 830 11595
rect 730 11515 830 11555
rect 730 11475 760 11515
rect 800 11475 830 11515
rect 730 11435 830 11475
rect 730 11395 760 11435
rect 800 11395 830 11435
rect 730 11355 830 11395
rect 730 11315 760 11355
rect 800 11315 830 11355
rect 730 11275 830 11315
rect 730 11235 760 11275
rect 800 11235 830 11275
rect 730 11195 830 11235
rect 730 11155 760 11195
rect 800 11155 830 11195
rect 730 11115 830 11155
rect 730 11075 760 11115
rect 800 11075 830 11115
rect 730 11035 830 11075
rect 730 10995 760 11035
rect 800 10995 830 11035
rect 730 10955 830 10995
rect 730 10915 760 10955
rect 800 10915 830 10955
rect 730 10875 830 10915
rect 730 10835 760 10875
rect 800 10835 830 10875
rect 730 10795 830 10835
rect 730 10755 760 10795
rect 800 10755 830 10795
rect 730 10715 830 10755
rect 730 10675 760 10715
rect 800 10675 830 10715
rect 730 10635 830 10675
rect 730 10595 760 10635
rect 800 10595 830 10635
rect 730 10555 830 10595
rect 730 10515 760 10555
rect 800 10515 830 10555
rect 730 10475 830 10515
rect 730 10435 760 10475
rect 800 10435 830 10475
rect 730 10395 830 10435
rect 730 10355 760 10395
rect 800 10355 830 10395
rect 730 10315 830 10355
rect 730 10275 760 10315
rect 800 10275 830 10315
rect 730 10245 830 10275
rect 845 12235 945 12270
rect 845 12195 875 12235
rect 915 12195 945 12235
rect 845 12155 945 12195
rect 845 12115 875 12155
rect 915 12115 945 12155
rect 845 12075 945 12115
rect 845 12035 875 12075
rect 915 12035 945 12075
rect 845 11995 945 12035
rect 845 11955 875 11995
rect 915 11955 945 11995
rect 845 11915 945 11955
rect 845 11875 875 11915
rect 915 11875 945 11915
rect 845 11835 945 11875
rect 845 11795 875 11835
rect 915 11795 945 11835
rect 845 11755 945 11795
rect 845 11715 875 11755
rect 915 11715 945 11755
rect 845 11675 945 11715
rect 845 11635 875 11675
rect 915 11635 945 11675
rect 845 11595 945 11635
rect 845 11555 875 11595
rect 915 11555 945 11595
rect 845 11515 945 11555
rect 845 11475 875 11515
rect 915 11475 945 11515
rect 845 11435 945 11475
rect 845 11395 875 11435
rect 915 11395 945 11435
rect 845 11355 945 11395
rect 845 11315 875 11355
rect 915 11315 945 11355
rect 845 11275 945 11315
rect 845 11235 875 11275
rect 915 11235 945 11275
rect 845 11195 945 11235
rect 845 11155 875 11195
rect 915 11155 945 11195
rect 845 11115 945 11155
rect 845 11075 875 11115
rect 915 11075 945 11115
rect 845 11035 945 11075
rect 845 10995 875 11035
rect 915 10995 945 11035
rect 845 10955 945 10995
rect 845 10915 875 10955
rect 915 10915 945 10955
rect 845 10875 945 10915
rect 845 10835 875 10875
rect 915 10835 945 10875
rect 845 10795 945 10835
rect 845 10755 875 10795
rect 915 10755 945 10795
rect 845 10715 945 10755
rect 845 10675 875 10715
rect 915 10675 945 10715
rect 845 10635 945 10675
rect 845 10595 875 10635
rect 915 10595 945 10635
rect 845 10555 945 10595
rect 845 10515 875 10555
rect 915 10515 945 10555
rect 845 10475 945 10515
rect 845 10435 875 10475
rect 915 10435 945 10475
rect 845 10395 945 10435
rect 845 10355 875 10395
rect 915 10355 945 10395
rect 845 10315 945 10355
rect 845 10275 875 10315
rect 915 10275 945 10315
rect 845 10245 945 10275
rect 960 12235 1060 12270
rect 960 12195 990 12235
rect 1030 12195 1060 12235
rect 960 12155 1060 12195
rect 960 12115 990 12155
rect 1030 12115 1060 12155
rect 960 12075 1060 12115
rect 960 12035 990 12075
rect 1030 12035 1060 12075
rect 960 11995 1060 12035
rect 960 11955 990 11995
rect 1030 11955 1060 11995
rect 960 11915 1060 11955
rect 960 11875 990 11915
rect 1030 11875 1060 11915
rect 960 11835 1060 11875
rect 960 11795 990 11835
rect 1030 11795 1060 11835
rect 960 11755 1060 11795
rect 960 11715 990 11755
rect 1030 11715 1060 11755
rect 960 11675 1060 11715
rect 960 11635 990 11675
rect 1030 11635 1060 11675
rect 960 11595 1060 11635
rect 960 11555 990 11595
rect 1030 11555 1060 11595
rect 960 11515 1060 11555
rect 960 11475 990 11515
rect 1030 11475 1060 11515
rect 960 11435 1060 11475
rect 960 11395 990 11435
rect 1030 11395 1060 11435
rect 960 11355 1060 11395
rect 960 11315 990 11355
rect 1030 11315 1060 11355
rect 960 11275 1060 11315
rect 960 11235 990 11275
rect 1030 11235 1060 11275
rect 960 11195 1060 11235
rect 960 11155 990 11195
rect 1030 11155 1060 11195
rect 960 11115 1060 11155
rect 960 11075 990 11115
rect 1030 11075 1060 11115
rect 960 11035 1060 11075
rect 960 10995 990 11035
rect 1030 10995 1060 11035
rect 960 10955 1060 10995
rect 960 10915 990 10955
rect 1030 10915 1060 10955
rect 960 10875 1060 10915
rect 960 10835 990 10875
rect 1030 10835 1060 10875
rect 960 10795 1060 10835
rect 960 10755 990 10795
rect 1030 10755 1060 10795
rect 960 10715 1060 10755
rect 960 10675 990 10715
rect 1030 10675 1060 10715
rect 960 10635 1060 10675
rect 960 10595 990 10635
rect 1030 10595 1060 10635
rect 960 10555 1060 10595
rect 960 10515 990 10555
rect 1030 10515 1060 10555
rect 960 10475 1060 10515
rect 960 10435 990 10475
rect 1030 10435 1060 10475
rect 960 10395 1060 10435
rect 960 10355 990 10395
rect 1030 10355 1060 10395
rect 960 10315 1060 10355
rect 960 10275 990 10315
rect 1030 10275 1060 10315
rect 960 10245 1060 10275
rect 1075 12235 1175 12270
rect 1075 12195 1105 12235
rect 1145 12195 1175 12235
rect 1075 12155 1175 12195
rect 1075 12115 1105 12155
rect 1145 12115 1175 12155
rect 1075 12075 1175 12115
rect 1075 12035 1105 12075
rect 1145 12035 1175 12075
rect 1075 11995 1175 12035
rect 1075 11955 1105 11995
rect 1145 11955 1175 11995
rect 1075 11915 1175 11955
rect 1075 11875 1105 11915
rect 1145 11875 1175 11915
rect 1075 11835 1175 11875
rect 1075 11795 1105 11835
rect 1145 11795 1175 11835
rect 1075 11755 1175 11795
rect 1075 11715 1105 11755
rect 1145 11715 1175 11755
rect 1075 11675 1175 11715
rect 1075 11635 1105 11675
rect 1145 11635 1175 11675
rect 1075 11595 1175 11635
rect 1075 11555 1105 11595
rect 1145 11555 1175 11595
rect 1075 11515 1175 11555
rect 1075 11475 1105 11515
rect 1145 11475 1175 11515
rect 1075 11435 1175 11475
rect 1075 11395 1105 11435
rect 1145 11395 1175 11435
rect 1075 11355 1175 11395
rect 1075 11315 1105 11355
rect 1145 11315 1175 11355
rect 1075 11275 1175 11315
rect 1075 11235 1105 11275
rect 1145 11235 1175 11275
rect 1075 11195 1175 11235
rect 1075 11155 1105 11195
rect 1145 11155 1175 11195
rect 1075 11115 1175 11155
rect 1075 11075 1105 11115
rect 1145 11075 1175 11115
rect 1075 11035 1175 11075
rect 1075 10995 1105 11035
rect 1145 10995 1175 11035
rect 1075 10955 1175 10995
rect 1075 10915 1105 10955
rect 1145 10915 1175 10955
rect 1075 10875 1175 10915
rect 1075 10835 1105 10875
rect 1145 10835 1175 10875
rect 1075 10795 1175 10835
rect 1075 10755 1105 10795
rect 1145 10755 1175 10795
rect 1075 10715 1175 10755
rect 1075 10675 1105 10715
rect 1145 10675 1175 10715
rect 1075 10635 1175 10675
rect 1075 10595 1105 10635
rect 1145 10595 1175 10635
rect 1075 10555 1175 10595
rect 1075 10515 1105 10555
rect 1145 10515 1175 10555
rect 1075 10475 1175 10515
rect 1075 10435 1105 10475
rect 1145 10435 1175 10475
rect 1075 10395 1175 10435
rect 1075 10355 1105 10395
rect 1145 10355 1175 10395
rect 1075 10315 1175 10355
rect 1075 10275 1105 10315
rect 1145 10275 1175 10315
rect 1075 10245 1175 10275
rect 1190 12235 1290 12270
rect 1190 12195 1220 12235
rect 1260 12195 1290 12235
rect 1190 12155 1290 12195
rect 1190 12115 1220 12155
rect 1260 12115 1290 12155
rect 1190 12075 1290 12115
rect 1190 12035 1220 12075
rect 1260 12035 1290 12075
rect 1190 11995 1290 12035
rect 1190 11955 1220 11995
rect 1260 11955 1290 11995
rect 1190 11915 1290 11955
rect 1190 11875 1220 11915
rect 1260 11875 1290 11915
rect 1190 11835 1290 11875
rect 1190 11795 1220 11835
rect 1260 11795 1290 11835
rect 1190 11755 1290 11795
rect 1190 11715 1220 11755
rect 1260 11715 1290 11755
rect 1190 11675 1290 11715
rect 1190 11635 1220 11675
rect 1260 11635 1290 11675
rect 1190 11595 1290 11635
rect 1190 11555 1220 11595
rect 1260 11555 1290 11595
rect 1190 11515 1290 11555
rect 1190 11475 1220 11515
rect 1260 11475 1290 11515
rect 1190 11435 1290 11475
rect 1190 11395 1220 11435
rect 1260 11395 1290 11435
rect 1190 11355 1290 11395
rect 1190 11315 1220 11355
rect 1260 11315 1290 11355
rect 1190 11275 1290 11315
rect 1190 11235 1220 11275
rect 1260 11235 1290 11275
rect 1190 11195 1290 11235
rect 1190 11155 1220 11195
rect 1260 11155 1290 11195
rect 1190 11115 1290 11155
rect 1190 11075 1220 11115
rect 1260 11075 1290 11115
rect 1190 11035 1290 11075
rect 1190 10995 1220 11035
rect 1260 10995 1290 11035
rect 1190 10955 1290 10995
rect 1190 10915 1220 10955
rect 1260 10915 1290 10955
rect 1190 10875 1290 10915
rect 1190 10835 1220 10875
rect 1260 10835 1290 10875
rect 1190 10795 1290 10835
rect 1190 10755 1220 10795
rect 1260 10755 1290 10795
rect 1190 10715 1290 10755
rect 1190 10675 1220 10715
rect 1260 10675 1290 10715
rect 1190 10635 1290 10675
rect 1190 10595 1220 10635
rect 1260 10595 1290 10635
rect 1190 10555 1290 10595
rect 1190 10515 1220 10555
rect 1260 10515 1290 10555
rect 1190 10475 1290 10515
rect 1190 10435 1220 10475
rect 1260 10435 1290 10475
rect 1190 10395 1290 10435
rect 1190 10355 1220 10395
rect 1260 10355 1290 10395
rect 1190 10315 1290 10355
rect 1190 10275 1220 10315
rect 1260 10275 1290 10315
rect 1190 10245 1290 10275
rect 1305 12235 1405 12270
rect 1305 12195 1335 12235
rect 1375 12195 1405 12235
rect 1305 12155 1405 12195
rect 1305 12115 1335 12155
rect 1375 12115 1405 12155
rect 1305 12075 1405 12115
rect 1305 12035 1335 12075
rect 1375 12035 1405 12075
rect 1305 11995 1405 12035
rect 1305 11955 1335 11995
rect 1375 11955 1405 11995
rect 1305 11915 1405 11955
rect 1305 11875 1335 11915
rect 1375 11875 1405 11915
rect 1305 11835 1405 11875
rect 1305 11795 1335 11835
rect 1375 11795 1405 11835
rect 1305 11755 1405 11795
rect 1305 11715 1335 11755
rect 1375 11715 1405 11755
rect 1305 11675 1405 11715
rect 1305 11635 1335 11675
rect 1375 11635 1405 11675
rect 1305 11595 1405 11635
rect 1305 11555 1335 11595
rect 1375 11555 1405 11595
rect 1305 11515 1405 11555
rect 1305 11475 1335 11515
rect 1375 11475 1405 11515
rect 1305 11435 1405 11475
rect 1305 11395 1335 11435
rect 1375 11395 1405 11435
rect 1305 11355 1405 11395
rect 1305 11315 1335 11355
rect 1375 11315 1405 11355
rect 1305 11275 1405 11315
rect 1305 11235 1335 11275
rect 1375 11235 1405 11275
rect 1305 11195 1405 11235
rect 1305 11155 1335 11195
rect 1375 11155 1405 11195
rect 1305 11115 1405 11155
rect 1305 11075 1335 11115
rect 1375 11075 1405 11115
rect 1305 11035 1405 11075
rect 1305 10995 1335 11035
rect 1375 10995 1405 11035
rect 1305 10955 1405 10995
rect 1305 10915 1335 10955
rect 1375 10915 1405 10955
rect 1305 10875 1405 10915
rect 1305 10835 1335 10875
rect 1375 10835 1405 10875
rect 1305 10795 1405 10835
rect 1305 10755 1335 10795
rect 1375 10755 1405 10795
rect 1305 10715 1405 10755
rect 1305 10675 1335 10715
rect 1375 10675 1405 10715
rect 1305 10635 1405 10675
rect 1305 10595 1335 10635
rect 1375 10595 1405 10635
rect 1305 10555 1405 10595
rect 1305 10515 1335 10555
rect 1375 10515 1405 10555
rect 1305 10475 1405 10515
rect 1305 10435 1335 10475
rect 1375 10435 1405 10475
rect 1305 10395 1405 10435
rect 1305 10355 1335 10395
rect 1375 10355 1405 10395
rect 1305 10315 1405 10355
rect 1305 10275 1335 10315
rect 1375 10275 1405 10315
rect 1305 10245 1405 10275
rect 1420 12235 1520 12270
rect 1420 12195 1450 12235
rect 1490 12195 1520 12235
rect 1420 12155 1520 12195
rect 1420 12115 1450 12155
rect 1490 12115 1520 12155
rect 1420 12075 1520 12115
rect 1420 12035 1450 12075
rect 1490 12035 1520 12075
rect 1420 11995 1520 12035
rect 1420 11955 1450 11995
rect 1490 11955 1520 11995
rect 1420 11915 1520 11955
rect 1420 11875 1450 11915
rect 1490 11875 1520 11915
rect 1420 11835 1520 11875
rect 1420 11795 1450 11835
rect 1490 11795 1520 11835
rect 1420 11755 1520 11795
rect 1420 11715 1450 11755
rect 1490 11715 1520 11755
rect 1420 11675 1520 11715
rect 1420 11635 1450 11675
rect 1490 11635 1520 11675
rect 1420 11595 1520 11635
rect 1420 11555 1450 11595
rect 1490 11555 1520 11595
rect 1420 11515 1520 11555
rect 1420 11475 1450 11515
rect 1490 11475 1520 11515
rect 1420 11435 1520 11475
rect 1420 11395 1450 11435
rect 1490 11395 1520 11435
rect 1420 11355 1520 11395
rect 1420 11315 1450 11355
rect 1490 11315 1520 11355
rect 1420 11275 1520 11315
rect 1420 11235 1450 11275
rect 1490 11235 1520 11275
rect 1420 11195 1520 11235
rect 1420 11155 1450 11195
rect 1490 11155 1520 11195
rect 1420 11115 1520 11155
rect 1420 11075 1450 11115
rect 1490 11075 1520 11115
rect 1420 11035 1520 11075
rect 1420 10995 1450 11035
rect 1490 10995 1520 11035
rect 1420 10955 1520 10995
rect 1420 10915 1450 10955
rect 1490 10915 1520 10955
rect 1420 10875 1520 10915
rect 1420 10835 1450 10875
rect 1490 10835 1520 10875
rect 1420 10795 1520 10835
rect 1420 10755 1450 10795
rect 1490 10755 1520 10795
rect 1420 10715 1520 10755
rect 1420 10675 1450 10715
rect 1490 10675 1520 10715
rect 1420 10635 1520 10675
rect 1420 10595 1450 10635
rect 1490 10595 1520 10635
rect 1420 10555 1520 10595
rect 1420 10515 1450 10555
rect 1490 10515 1520 10555
rect 1420 10475 1520 10515
rect 1420 10435 1450 10475
rect 1490 10435 1520 10475
rect 1420 10395 1520 10435
rect 1420 10355 1450 10395
rect 1490 10355 1520 10395
rect 1420 10315 1520 10355
rect 1420 10275 1450 10315
rect 1490 10275 1520 10315
rect 1420 10245 1520 10275
rect 1535 12235 1635 12270
rect 1535 12195 1565 12235
rect 1605 12195 1635 12235
rect 1535 12155 1635 12195
rect 1535 12115 1565 12155
rect 1605 12115 1635 12155
rect 1535 12075 1635 12115
rect 1535 12035 1565 12075
rect 1605 12035 1635 12075
rect 1535 11995 1635 12035
rect 1535 11955 1565 11995
rect 1605 11955 1635 11995
rect 1535 11915 1635 11955
rect 1535 11875 1565 11915
rect 1605 11875 1635 11915
rect 1535 11835 1635 11875
rect 1535 11795 1565 11835
rect 1605 11795 1635 11835
rect 1535 11755 1635 11795
rect 1535 11715 1565 11755
rect 1605 11715 1635 11755
rect 1535 11675 1635 11715
rect 1535 11635 1565 11675
rect 1605 11635 1635 11675
rect 1535 11595 1635 11635
rect 1535 11555 1565 11595
rect 1605 11555 1635 11595
rect 1535 11515 1635 11555
rect 1535 11475 1565 11515
rect 1605 11475 1635 11515
rect 1535 11435 1635 11475
rect 1535 11395 1565 11435
rect 1605 11395 1635 11435
rect 1535 11355 1635 11395
rect 1535 11315 1565 11355
rect 1605 11315 1635 11355
rect 1535 11275 1635 11315
rect 1535 11235 1565 11275
rect 1605 11235 1635 11275
rect 1535 11195 1635 11235
rect 1535 11155 1565 11195
rect 1605 11155 1635 11195
rect 1535 11115 1635 11155
rect 1535 11075 1565 11115
rect 1605 11075 1635 11115
rect 1535 11035 1635 11075
rect 1535 10995 1565 11035
rect 1605 10995 1635 11035
rect 1535 10955 1635 10995
rect 1535 10915 1565 10955
rect 1605 10915 1635 10955
rect 1535 10875 1635 10915
rect 1535 10835 1565 10875
rect 1605 10835 1635 10875
rect 1535 10795 1635 10835
rect 1535 10755 1565 10795
rect 1605 10755 1635 10795
rect 1535 10715 1635 10755
rect 1535 10675 1565 10715
rect 1605 10675 1635 10715
rect 1535 10635 1635 10675
rect 1535 10595 1565 10635
rect 1605 10595 1635 10635
rect 1535 10555 1635 10595
rect 1535 10515 1565 10555
rect 1605 10515 1635 10555
rect 1535 10475 1635 10515
rect 1535 10435 1565 10475
rect 1605 10435 1635 10475
rect 1535 10395 1635 10435
rect 1535 10355 1565 10395
rect 1605 10355 1635 10395
rect 1535 10315 1635 10355
rect 1535 10275 1565 10315
rect 1605 10275 1635 10315
rect 1535 10245 1635 10275
rect 1650 12235 1750 12270
rect 1650 12195 1680 12235
rect 1720 12195 1750 12235
rect 1650 12155 1750 12195
rect 1650 12115 1680 12155
rect 1720 12115 1750 12155
rect 1650 12075 1750 12115
rect 1650 12035 1680 12075
rect 1720 12035 1750 12075
rect 1650 11995 1750 12035
rect 1650 11955 1680 11995
rect 1720 11955 1750 11995
rect 1650 11915 1750 11955
rect 1650 11875 1680 11915
rect 1720 11875 1750 11915
rect 1650 11835 1750 11875
rect 1650 11795 1680 11835
rect 1720 11795 1750 11835
rect 1650 11755 1750 11795
rect 1650 11715 1680 11755
rect 1720 11715 1750 11755
rect 1650 11675 1750 11715
rect 1650 11635 1680 11675
rect 1720 11635 1750 11675
rect 1650 11595 1750 11635
rect 1650 11555 1680 11595
rect 1720 11555 1750 11595
rect 1650 11515 1750 11555
rect 1650 11475 1680 11515
rect 1720 11475 1750 11515
rect 1650 11435 1750 11475
rect 1650 11395 1680 11435
rect 1720 11395 1750 11435
rect 1650 11355 1750 11395
rect 1650 11315 1680 11355
rect 1720 11315 1750 11355
rect 1650 11275 1750 11315
rect 1650 11235 1680 11275
rect 1720 11235 1750 11275
rect 1650 11195 1750 11235
rect 1650 11155 1680 11195
rect 1720 11155 1750 11195
rect 1650 11115 1750 11155
rect 1650 11075 1680 11115
rect 1720 11075 1750 11115
rect 1650 11035 1750 11075
rect 1650 10995 1680 11035
rect 1720 10995 1750 11035
rect 1650 10955 1750 10995
rect 1650 10915 1680 10955
rect 1720 10915 1750 10955
rect 1650 10875 1750 10915
rect 1650 10835 1680 10875
rect 1720 10835 1750 10875
rect 1650 10795 1750 10835
rect 1650 10755 1680 10795
rect 1720 10755 1750 10795
rect 1650 10715 1750 10755
rect 1650 10675 1680 10715
rect 1720 10675 1750 10715
rect 1650 10635 1750 10675
rect 1650 10595 1680 10635
rect 1720 10595 1750 10635
rect 1650 10555 1750 10595
rect 1650 10515 1680 10555
rect 1720 10515 1750 10555
rect 1650 10475 1750 10515
rect 1650 10435 1680 10475
rect 1720 10435 1750 10475
rect 1650 10395 1750 10435
rect 1650 10355 1680 10395
rect 1720 10355 1750 10395
rect 1650 10315 1750 10355
rect 1650 10275 1680 10315
rect 1720 10275 1750 10315
rect 1650 10245 1750 10275
rect 1765 12235 1865 12270
rect 1765 12195 1795 12235
rect 1835 12195 1865 12235
rect 1765 12155 1865 12195
rect 1765 12115 1795 12155
rect 1835 12115 1865 12155
rect 1765 12075 1865 12115
rect 1765 12035 1795 12075
rect 1835 12035 1865 12075
rect 1765 11995 1865 12035
rect 1765 11955 1795 11995
rect 1835 11955 1865 11995
rect 1765 11915 1865 11955
rect 1765 11875 1795 11915
rect 1835 11875 1865 11915
rect 1765 11835 1865 11875
rect 1765 11795 1795 11835
rect 1835 11795 1865 11835
rect 1765 11755 1865 11795
rect 1765 11715 1795 11755
rect 1835 11715 1865 11755
rect 1765 11675 1865 11715
rect 1765 11635 1795 11675
rect 1835 11635 1865 11675
rect 1765 11595 1865 11635
rect 1765 11555 1795 11595
rect 1835 11555 1865 11595
rect 1765 11515 1865 11555
rect 1765 11475 1795 11515
rect 1835 11475 1865 11515
rect 1765 11435 1865 11475
rect 1765 11395 1795 11435
rect 1835 11395 1865 11435
rect 1765 11355 1865 11395
rect 1765 11315 1795 11355
rect 1835 11315 1865 11355
rect 1765 11275 1865 11315
rect 1765 11235 1795 11275
rect 1835 11235 1865 11275
rect 1765 11195 1865 11235
rect 1765 11155 1795 11195
rect 1835 11155 1865 11195
rect 1765 11115 1865 11155
rect 1765 11075 1795 11115
rect 1835 11075 1865 11115
rect 1765 11035 1865 11075
rect 1765 10995 1795 11035
rect 1835 10995 1865 11035
rect 1765 10955 1865 10995
rect 1765 10915 1795 10955
rect 1835 10915 1865 10955
rect 1765 10875 1865 10915
rect 1765 10835 1795 10875
rect 1835 10835 1865 10875
rect 1765 10795 1865 10835
rect 1765 10755 1795 10795
rect 1835 10755 1865 10795
rect 1765 10715 1865 10755
rect 1765 10675 1795 10715
rect 1835 10675 1865 10715
rect 1765 10635 1865 10675
rect 1765 10595 1795 10635
rect 1835 10595 1865 10635
rect 1765 10555 1865 10595
rect 1765 10515 1795 10555
rect 1835 10515 1865 10555
rect 1765 10475 1865 10515
rect 1765 10435 1795 10475
rect 1835 10435 1865 10475
rect 1765 10395 1865 10435
rect 1765 10355 1795 10395
rect 1835 10355 1865 10395
rect 1765 10315 1865 10355
rect 1765 10275 1795 10315
rect 1835 10275 1865 10315
rect 1765 10245 1865 10275
rect 1880 12235 1980 12270
rect 1880 12195 1910 12235
rect 1950 12195 1980 12235
rect 1880 12155 1980 12195
rect 1880 12115 1910 12155
rect 1950 12115 1980 12155
rect 1880 12075 1980 12115
rect 1880 12035 1910 12075
rect 1950 12035 1980 12075
rect 1880 11995 1980 12035
rect 1880 11955 1910 11995
rect 1950 11955 1980 11995
rect 1880 11915 1980 11955
rect 1880 11875 1910 11915
rect 1950 11875 1980 11915
rect 1880 11835 1980 11875
rect 1880 11795 1910 11835
rect 1950 11795 1980 11835
rect 1880 11755 1980 11795
rect 1880 11715 1910 11755
rect 1950 11715 1980 11755
rect 1880 11675 1980 11715
rect 1880 11635 1910 11675
rect 1950 11635 1980 11675
rect 1880 11595 1980 11635
rect 1880 11555 1910 11595
rect 1950 11555 1980 11595
rect 1880 11515 1980 11555
rect 1880 11475 1910 11515
rect 1950 11475 1980 11515
rect 1880 11435 1980 11475
rect 1880 11395 1910 11435
rect 1950 11395 1980 11435
rect 1880 11355 1980 11395
rect 1880 11315 1910 11355
rect 1950 11315 1980 11355
rect 1880 11275 1980 11315
rect 1880 11235 1910 11275
rect 1950 11235 1980 11275
rect 1880 11195 1980 11235
rect 1880 11155 1910 11195
rect 1950 11155 1980 11195
rect 1880 11115 1980 11155
rect 1880 11075 1910 11115
rect 1950 11075 1980 11115
rect 1880 11035 1980 11075
rect 1880 10995 1910 11035
rect 1950 10995 1980 11035
rect 1880 10955 1980 10995
rect 1880 10915 1910 10955
rect 1950 10915 1980 10955
rect 1880 10875 1980 10915
rect 1880 10835 1910 10875
rect 1950 10835 1980 10875
rect 1880 10795 1980 10835
rect 1880 10755 1910 10795
rect 1950 10755 1980 10795
rect 1880 10715 1980 10755
rect 1880 10675 1910 10715
rect 1950 10675 1980 10715
rect 1880 10635 1980 10675
rect 1880 10595 1910 10635
rect 1950 10595 1980 10635
rect 1880 10555 1980 10595
rect 1880 10515 1910 10555
rect 1950 10515 1980 10555
rect 1880 10475 1980 10515
rect 1880 10435 1910 10475
rect 1950 10435 1980 10475
rect 1880 10395 1980 10435
rect 1880 10355 1910 10395
rect 1950 10355 1980 10395
rect 1880 10315 1980 10355
rect 1880 10275 1910 10315
rect 1950 10275 1980 10315
rect 1880 10245 1980 10275
rect 1995 12235 2095 12270
rect 1995 12195 2025 12235
rect 2065 12195 2095 12235
rect 1995 12155 2095 12195
rect 1995 12115 2025 12155
rect 2065 12115 2095 12155
rect 1995 12075 2095 12115
rect 1995 12035 2025 12075
rect 2065 12035 2095 12075
rect 1995 11995 2095 12035
rect 1995 11955 2025 11995
rect 2065 11955 2095 11995
rect 1995 11915 2095 11955
rect 1995 11875 2025 11915
rect 2065 11875 2095 11915
rect 1995 11835 2095 11875
rect 1995 11795 2025 11835
rect 2065 11795 2095 11835
rect 1995 11755 2095 11795
rect 1995 11715 2025 11755
rect 2065 11715 2095 11755
rect 1995 11675 2095 11715
rect 1995 11635 2025 11675
rect 2065 11635 2095 11675
rect 1995 11595 2095 11635
rect 1995 11555 2025 11595
rect 2065 11555 2095 11595
rect 1995 11515 2095 11555
rect 1995 11475 2025 11515
rect 2065 11475 2095 11515
rect 1995 11435 2095 11475
rect 1995 11395 2025 11435
rect 2065 11395 2095 11435
rect 1995 11355 2095 11395
rect 1995 11315 2025 11355
rect 2065 11315 2095 11355
rect 1995 11275 2095 11315
rect 1995 11235 2025 11275
rect 2065 11235 2095 11275
rect 1995 11195 2095 11235
rect 1995 11155 2025 11195
rect 2065 11155 2095 11195
rect 1995 11115 2095 11155
rect 1995 11075 2025 11115
rect 2065 11075 2095 11115
rect 1995 11035 2095 11075
rect 1995 10995 2025 11035
rect 2065 10995 2095 11035
rect 1995 10955 2095 10995
rect 1995 10915 2025 10955
rect 2065 10915 2095 10955
rect 1995 10875 2095 10915
rect 1995 10835 2025 10875
rect 2065 10835 2095 10875
rect 1995 10795 2095 10835
rect 1995 10755 2025 10795
rect 2065 10755 2095 10795
rect 1995 10715 2095 10755
rect 1995 10675 2025 10715
rect 2065 10675 2095 10715
rect 1995 10635 2095 10675
rect 1995 10595 2025 10635
rect 2065 10595 2095 10635
rect 1995 10555 2095 10595
rect 1995 10515 2025 10555
rect 2065 10515 2095 10555
rect 1995 10475 2095 10515
rect 1995 10435 2025 10475
rect 2065 10435 2095 10475
rect 1995 10395 2095 10435
rect 1995 10355 2025 10395
rect 2065 10355 2095 10395
rect 1995 10315 2095 10355
rect 1995 10275 2025 10315
rect 2065 10275 2095 10315
rect 1995 10245 2095 10275
rect 2110 12235 2210 12270
rect 2110 12195 2140 12235
rect 2180 12195 2210 12235
rect 2110 12155 2210 12195
rect 2110 12115 2140 12155
rect 2180 12115 2210 12155
rect 2110 12075 2210 12115
rect 2110 12035 2140 12075
rect 2180 12035 2210 12075
rect 2110 11995 2210 12035
rect 2110 11955 2140 11995
rect 2180 11955 2210 11995
rect 2110 11915 2210 11955
rect 2110 11875 2140 11915
rect 2180 11875 2210 11915
rect 2110 11835 2210 11875
rect 2110 11795 2140 11835
rect 2180 11795 2210 11835
rect 2110 11755 2210 11795
rect 2110 11715 2140 11755
rect 2180 11715 2210 11755
rect 2110 11675 2210 11715
rect 2110 11635 2140 11675
rect 2180 11635 2210 11675
rect 2110 11595 2210 11635
rect 2110 11555 2140 11595
rect 2180 11555 2210 11595
rect 2110 11515 2210 11555
rect 2110 11475 2140 11515
rect 2180 11475 2210 11515
rect 2110 11435 2210 11475
rect 2110 11395 2140 11435
rect 2180 11395 2210 11435
rect 2110 11355 2210 11395
rect 2110 11315 2140 11355
rect 2180 11315 2210 11355
rect 2110 11275 2210 11315
rect 2110 11235 2140 11275
rect 2180 11235 2210 11275
rect 2110 11195 2210 11235
rect 2110 11155 2140 11195
rect 2180 11155 2210 11195
rect 2110 11115 2210 11155
rect 2110 11075 2140 11115
rect 2180 11075 2210 11115
rect 2110 11035 2210 11075
rect 2110 10995 2140 11035
rect 2180 10995 2210 11035
rect 2110 10955 2210 10995
rect 2110 10915 2140 10955
rect 2180 10915 2210 10955
rect 2110 10875 2210 10915
rect 2110 10835 2140 10875
rect 2180 10835 2210 10875
rect 2110 10795 2210 10835
rect 2110 10755 2140 10795
rect 2180 10755 2210 10795
rect 2110 10715 2210 10755
rect 2110 10675 2140 10715
rect 2180 10675 2210 10715
rect 2110 10635 2210 10675
rect 2110 10595 2140 10635
rect 2180 10595 2210 10635
rect 2110 10555 2210 10595
rect 2110 10515 2140 10555
rect 2180 10515 2210 10555
rect 2110 10475 2210 10515
rect 2110 10435 2140 10475
rect 2180 10435 2210 10475
rect 2110 10395 2210 10435
rect 2110 10355 2140 10395
rect 2180 10355 2210 10395
rect 2110 10315 2210 10355
rect 2110 10275 2140 10315
rect 2180 10275 2210 10315
rect 2110 10245 2210 10275
rect 2225 12235 2325 12270
rect 2225 12195 2255 12235
rect 2295 12195 2325 12235
rect 2225 12155 2325 12195
rect 2225 12115 2255 12155
rect 2295 12115 2325 12155
rect 2225 12075 2325 12115
rect 2225 12035 2255 12075
rect 2295 12035 2325 12075
rect 2225 11995 2325 12035
rect 2225 11955 2255 11995
rect 2295 11955 2325 11995
rect 2225 11915 2325 11955
rect 2225 11875 2255 11915
rect 2295 11875 2325 11915
rect 2225 11835 2325 11875
rect 2225 11795 2255 11835
rect 2295 11795 2325 11835
rect 2225 11755 2325 11795
rect 2225 11715 2255 11755
rect 2295 11715 2325 11755
rect 2225 11675 2325 11715
rect 2225 11635 2255 11675
rect 2295 11635 2325 11675
rect 2225 11595 2325 11635
rect 2225 11555 2255 11595
rect 2295 11555 2325 11595
rect 2225 11515 2325 11555
rect 2225 11475 2255 11515
rect 2295 11475 2325 11515
rect 2225 11435 2325 11475
rect 2225 11395 2255 11435
rect 2295 11395 2325 11435
rect 2225 11355 2325 11395
rect 2225 11315 2255 11355
rect 2295 11315 2325 11355
rect 2225 11275 2325 11315
rect 2225 11235 2255 11275
rect 2295 11235 2325 11275
rect 2225 11195 2325 11235
rect 2225 11155 2255 11195
rect 2295 11155 2325 11195
rect 2225 11115 2325 11155
rect 2225 11075 2255 11115
rect 2295 11075 2325 11115
rect 2225 11035 2325 11075
rect 2225 10995 2255 11035
rect 2295 10995 2325 11035
rect 2225 10955 2325 10995
rect 2225 10915 2255 10955
rect 2295 10915 2325 10955
rect 2225 10875 2325 10915
rect 2225 10835 2255 10875
rect 2295 10835 2325 10875
rect 2225 10795 2325 10835
rect 2225 10755 2255 10795
rect 2295 10755 2325 10795
rect 2225 10715 2325 10755
rect 2225 10675 2255 10715
rect 2295 10675 2325 10715
rect 2225 10635 2325 10675
rect 2225 10595 2255 10635
rect 2295 10595 2325 10635
rect 2225 10555 2325 10595
rect 2225 10515 2255 10555
rect 2295 10515 2325 10555
rect 2225 10475 2325 10515
rect 2225 10435 2255 10475
rect 2295 10435 2325 10475
rect 2225 10395 2325 10435
rect 2225 10355 2255 10395
rect 2295 10355 2325 10395
rect 2225 10315 2325 10355
rect 2225 10275 2255 10315
rect 2295 10275 2325 10315
rect 2225 10245 2325 10275
rect 2340 12235 2440 12270
rect 2340 12195 2370 12235
rect 2410 12195 2440 12235
rect 2340 12155 2440 12195
rect 2340 12115 2370 12155
rect 2410 12115 2440 12155
rect 2340 12075 2440 12115
rect 2340 12035 2370 12075
rect 2410 12035 2440 12075
rect 2340 11995 2440 12035
rect 2340 11955 2370 11995
rect 2410 11955 2440 11995
rect 2340 11915 2440 11955
rect 2340 11875 2370 11915
rect 2410 11875 2440 11915
rect 2340 11835 2440 11875
rect 2340 11795 2370 11835
rect 2410 11795 2440 11835
rect 2340 11755 2440 11795
rect 2340 11715 2370 11755
rect 2410 11715 2440 11755
rect 2340 11675 2440 11715
rect 2340 11635 2370 11675
rect 2410 11635 2440 11675
rect 2340 11595 2440 11635
rect 2340 11555 2370 11595
rect 2410 11555 2440 11595
rect 2340 11515 2440 11555
rect 2340 11475 2370 11515
rect 2410 11475 2440 11515
rect 2340 11435 2440 11475
rect 2340 11395 2370 11435
rect 2410 11395 2440 11435
rect 2340 11355 2440 11395
rect 2340 11315 2370 11355
rect 2410 11315 2440 11355
rect 2340 11275 2440 11315
rect 2340 11235 2370 11275
rect 2410 11235 2440 11275
rect 2340 11195 2440 11235
rect 2340 11155 2370 11195
rect 2410 11155 2440 11195
rect 2340 11115 2440 11155
rect 2340 11075 2370 11115
rect 2410 11075 2440 11115
rect 2340 11035 2440 11075
rect 2340 10995 2370 11035
rect 2410 10995 2440 11035
rect 2340 10955 2440 10995
rect 2340 10915 2370 10955
rect 2410 10915 2440 10955
rect 2340 10875 2440 10915
rect 2340 10835 2370 10875
rect 2410 10835 2440 10875
rect 2340 10795 2440 10835
rect 2340 10755 2370 10795
rect 2410 10755 2440 10795
rect 2340 10715 2440 10755
rect 2340 10675 2370 10715
rect 2410 10675 2440 10715
rect 2340 10635 2440 10675
rect 2340 10595 2370 10635
rect 2410 10595 2440 10635
rect 2340 10555 2440 10595
rect 2340 10515 2370 10555
rect 2410 10515 2440 10555
rect 2340 10475 2440 10515
rect 2340 10435 2370 10475
rect 2410 10435 2440 10475
rect 2340 10395 2440 10435
rect 2340 10355 2370 10395
rect 2410 10355 2440 10395
rect 2340 10315 2440 10355
rect 2340 10275 2370 10315
rect 2410 10275 2440 10315
rect 2340 10245 2440 10275
rect 2455 12235 2555 12270
rect 2455 12195 2485 12235
rect 2525 12195 2555 12235
rect 2455 12155 2555 12195
rect 2455 12115 2485 12155
rect 2525 12115 2555 12155
rect 2455 12075 2555 12115
rect 2455 12035 2485 12075
rect 2525 12035 2555 12075
rect 2455 11995 2555 12035
rect 2455 11955 2485 11995
rect 2525 11955 2555 11995
rect 2455 11915 2555 11955
rect 2455 11875 2485 11915
rect 2525 11875 2555 11915
rect 2455 11835 2555 11875
rect 2455 11795 2485 11835
rect 2525 11795 2555 11835
rect 2455 11755 2555 11795
rect 2455 11715 2485 11755
rect 2525 11715 2555 11755
rect 2455 11675 2555 11715
rect 2455 11635 2485 11675
rect 2525 11635 2555 11675
rect 2455 11595 2555 11635
rect 2455 11555 2485 11595
rect 2525 11555 2555 11595
rect 2455 11515 2555 11555
rect 2455 11475 2485 11515
rect 2525 11475 2555 11515
rect 2455 11435 2555 11475
rect 2455 11395 2485 11435
rect 2525 11395 2555 11435
rect 2455 11355 2555 11395
rect 2455 11315 2485 11355
rect 2525 11315 2555 11355
rect 2455 11275 2555 11315
rect 2455 11235 2485 11275
rect 2525 11235 2555 11275
rect 2455 11195 2555 11235
rect 2455 11155 2485 11195
rect 2525 11155 2555 11195
rect 2455 11115 2555 11155
rect 2455 11075 2485 11115
rect 2525 11075 2555 11115
rect 2455 11035 2555 11075
rect 2455 10995 2485 11035
rect 2525 10995 2555 11035
rect 2455 10955 2555 10995
rect 2455 10915 2485 10955
rect 2525 10915 2555 10955
rect 2455 10875 2555 10915
rect 2455 10835 2485 10875
rect 2525 10835 2555 10875
rect 2455 10795 2555 10835
rect 2455 10755 2485 10795
rect 2525 10755 2555 10795
rect 2455 10715 2555 10755
rect 2455 10675 2485 10715
rect 2525 10675 2555 10715
rect 2455 10635 2555 10675
rect 2455 10595 2485 10635
rect 2525 10595 2555 10635
rect 2455 10555 2555 10595
rect 2455 10515 2485 10555
rect 2525 10515 2555 10555
rect 2455 10475 2555 10515
rect 2455 10435 2485 10475
rect 2525 10435 2555 10475
rect 2455 10395 2555 10435
rect 2455 10355 2485 10395
rect 2525 10355 2555 10395
rect 2455 10315 2555 10355
rect 2455 10275 2485 10315
rect 2525 10275 2555 10315
rect 2455 10245 2555 10275
<< pdiffc >>
rect -390 12195 -350 12235
rect -390 12115 -350 12155
rect -390 12035 -350 12075
rect -390 11955 -350 11995
rect -390 11875 -350 11915
rect -390 11795 -350 11835
rect -390 11715 -350 11755
rect -390 11635 -350 11675
rect -390 11555 -350 11595
rect -390 11475 -350 11515
rect -390 11395 -350 11435
rect -390 11315 -350 11355
rect -390 11235 -350 11275
rect -390 11155 -350 11195
rect -390 11075 -350 11115
rect -390 10995 -350 11035
rect -390 10915 -350 10955
rect -390 10835 -350 10875
rect -390 10755 -350 10795
rect -390 10675 -350 10715
rect -390 10595 -350 10635
rect -390 10515 -350 10555
rect -390 10435 -350 10475
rect -390 10355 -350 10395
rect -390 10275 -350 10315
rect -275 12195 -235 12235
rect -275 12115 -235 12155
rect -275 12035 -235 12075
rect -275 11955 -235 11995
rect -275 11875 -235 11915
rect -275 11795 -235 11835
rect -275 11715 -235 11755
rect -275 11635 -235 11675
rect -275 11555 -235 11595
rect -275 11475 -235 11515
rect -275 11395 -235 11435
rect -275 11315 -235 11355
rect -275 11235 -235 11275
rect -275 11155 -235 11195
rect -275 11075 -235 11115
rect -275 10995 -235 11035
rect -275 10915 -235 10955
rect -275 10835 -235 10875
rect -275 10755 -235 10795
rect -275 10675 -235 10715
rect -275 10595 -235 10635
rect -275 10515 -235 10555
rect -275 10435 -235 10475
rect -275 10355 -235 10395
rect -275 10275 -235 10315
rect -160 12195 -120 12235
rect -160 12115 -120 12155
rect -160 12035 -120 12075
rect -160 11955 -120 11995
rect -160 11875 -120 11915
rect -160 11795 -120 11835
rect -160 11715 -120 11755
rect -160 11635 -120 11675
rect -160 11555 -120 11595
rect -160 11475 -120 11515
rect -160 11395 -120 11435
rect -160 11315 -120 11355
rect -160 11235 -120 11275
rect -160 11155 -120 11195
rect -160 11075 -120 11115
rect -160 10995 -120 11035
rect -160 10915 -120 10955
rect -160 10835 -120 10875
rect -160 10755 -120 10795
rect -160 10675 -120 10715
rect -160 10595 -120 10635
rect -160 10515 -120 10555
rect -160 10435 -120 10475
rect -160 10355 -120 10395
rect -160 10275 -120 10315
rect -45 12195 -5 12235
rect -45 12115 -5 12155
rect -45 12035 -5 12075
rect -45 11955 -5 11995
rect -45 11875 -5 11915
rect -45 11795 -5 11835
rect -45 11715 -5 11755
rect -45 11635 -5 11675
rect -45 11555 -5 11595
rect -45 11475 -5 11515
rect -45 11395 -5 11435
rect -45 11315 -5 11355
rect -45 11235 -5 11275
rect -45 11155 -5 11195
rect -45 11075 -5 11115
rect -45 10995 -5 11035
rect -45 10915 -5 10955
rect -45 10835 -5 10875
rect -45 10755 -5 10795
rect -45 10675 -5 10715
rect -45 10595 -5 10635
rect -45 10515 -5 10555
rect -45 10435 -5 10475
rect -45 10355 -5 10395
rect -45 10275 -5 10315
rect 70 12195 110 12235
rect 70 12115 110 12155
rect 70 12035 110 12075
rect 70 11955 110 11995
rect 70 11875 110 11915
rect 70 11795 110 11835
rect 70 11715 110 11755
rect 70 11635 110 11675
rect 70 11555 110 11595
rect 70 11475 110 11515
rect 70 11395 110 11435
rect 70 11315 110 11355
rect 70 11235 110 11275
rect 70 11155 110 11195
rect 70 11075 110 11115
rect 70 10995 110 11035
rect 70 10915 110 10955
rect 70 10835 110 10875
rect 70 10755 110 10795
rect 70 10675 110 10715
rect 70 10595 110 10635
rect 70 10515 110 10555
rect 70 10435 110 10475
rect 70 10355 110 10395
rect 70 10275 110 10315
rect 185 12195 225 12235
rect 185 12115 225 12155
rect 185 12035 225 12075
rect 185 11955 225 11995
rect 185 11875 225 11915
rect 185 11795 225 11835
rect 185 11715 225 11755
rect 185 11635 225 11675
rect 185 11555 225 11595
rect 185 11475 225 11515
rect 185 11395 225 11435
rect 185 11315 225 11355
rect 185 11235 225 11275
rect 185 11155 225 11195
rect 185 11075 225 11115
rect 185 10995 225 11035
rect 185 10915 225 10955
rect 185 10835 225 10875
rect 185 10755 225 10795
rect 185 10675 225 10715
rect 185 10595 225 10635
rect 185 10515 225 10555
rect 185 10435 225 10475
rect 185 10355 225 10395
rect 185 10275 225 10315
rect 300 12195 340 12235
rect 300 12115 340 12155
rect 300 12035 340 12075
rect 300 11955 340 11995
rect 300 11875 340 11915
rect 300 11795 340 11835
rect 300 11715 340 11755
rect 300 11635 340 11675
rect 300 11555 340 11595
rect 300 11475 340 11515
rect 300 11395 340 11435
rect 300 11315 340 11355
rect 300 11235 340 11275
rect 300 11155 340 11195
rect 300 11075 340 11115
rect 300 10995 340 11035
rect 300 10915 340 10955
rect 300 10835 340 10875
rect 300 10755 340 10795
rect 300 10675 340 10715
rect 300 10595 340 10635
rect 300 10515 340 10555
rect 300 10435 340 10475
rect 300 10355 340 10395
rect 300 10275 340 10315
rect 415 12195 455 12235
rect 415 12115 455 12155
rect 415 12035 455 12075
rect 415 11955 455 11995
rect 415 11875 455 11915
rect 415 11795 455 11835
rect 415 11715 455 11755
rect 415 11635 455 11675
rect 415 11555 455 11595
rect 415 11475 455 11515
rect 415 11395 455 11435
rect 415 11315 455 11355
rect 415 11235 455 11275
rect 415 11155 455 11195
rect 415 11075 455 11115
rect 415 10995 455 11035
rect 415 10915 455 10955
rect 415 10835 455 10875
rect 415 10755 455 10795
rect 415 10675 455 10715
rect 415 10595 455 10635
rect 415 10515 455 10555
rect 415 10435 455 10475
rect 415 10355 455 10395
rect 415 10275 455 10315
rect 530 12195 570 12235
rect 530 12115 570 12155
rect 530 12035 570 12075
rect 530 11955 570 11995
rect 530 11875 570 11915
rect 530 11795 570 11835
rect 530 11715 570 11755
rect 530 11635 570 11675
rect 530 11555 570 11595
rect 530 11475 570 11515
rect 530 11395 570 11435
rect 530 11315 570 11355
rect 530 11235 570 11275
rect 530 11155 570 11195
rect 530 11075 570 11115
rect 530 10995 570 11035
rect 530 10915 570 10955
rect 530 10835 570 10875
rect 530 10755 570 10795
rect 530 10675 570 10715
rect 530 10595 570 10635
rect 530 10515 570 10555
rect 530 10435 570 10475
rect 530 10355 570 10395
rect 530 10275 570 10315
rect 645 12195 685 12235
rect 645 12115 685 12155
rect 645 12035 685 12075
rect 645 11955 685 11995
rect 645 11875 685 11915
rect 645 11795 685 11835
rect 645 11715 685 11755
rect 645 11635 685 11675
rect 645 11555 685 11595
rect 645 11475 685 11515
rect 645 11395 685 11435
rect 645 11315 685 11355
rect 645 11235 685 11275
rect 645 11155 685 11195
rect 645 11075 685 11115
rect 645 10995 685 11035
rect 645 10915 685 10955
rect 645 10835 685 10875
rect 645 10755 685 10795
rect 645 10675 685 10715
rect 645 10595 685 10635
rect 645 10515 685 10555
rect 645 10435 685 10475
rect 645 10355 685 10395
rect 645 10275 685 10315
rect 760 12195 800 12235
rect 760 12115 800 12155
rect 760 12035 800 12075
rect 760 11955 800 11995
rect 760 11875 800 11915
rect 760 11795 800 11835
rect 760 11715 800 11755
rect 760 11635 800 11675
rect 760 11555 800 11595
rect 760 11475 800 11515
rect 760 11395 800 11435
rect 760 11315 800 11355
rect 760 11235 800 11275
rect 760 11155 800 11195
rect 760 11075 800 11115
rect 760 10995 800 11035
rect 760 10915 800 10955
rect 760 10835 800 10875
rect 760 10755 800 10795
rect 760 10675 800 10715
rect 760 10595 800 10635
rect 760 10515 800 10555
rect 760 10435 800 10475
rect 760 10355 800 10395
rect 760 10275 800 10315
rect 875 12195 915 12235
rect 875 12115 915 12155
rect 875 12035 915 12075
rect 875 11955 915 11995
rect 875 11875 915 11915
rect 875 11795 915 11835
rect 875 11715 915 11755
rect 875 11635 915 11675
rect 875 11555 915 11595
rect 875 11475 915 11515
rect 875 11395 915 11435
rect 875 11315 915 11355
rect 875 11235 915 11275
rect 875 11155 915 11195
rect 875 11075 915 11115
rect 875 10995 915 11035
rect 875 10915 915 10955
rect 875 10835 915 10875
rect 875 10755 915 10795
rect 875 10675 915 10715
rect 875 10595 915 10635
rect 875 10515 915 10555
rect 875 10435 915 10475
rect 875 10355 915 10395
rect 875 10275 915 10315
rect 990 12195 1030 12235
rect 990 12115 1030 12155
rect 990 12035 1030 12075
rect 990 11955 1030 11995
rect 990 11875 1030 11915
rect 990 11795 1030 11835
rect 990 11715 1030 11755
rect 990 11635 1030 11675
rect 990 11555 1030 11595
rect 990 11475 1030 11515
rect 990 11395 1030 11435
rect 990 11315 1030 11355
rect 990 11235 1030 11275
rect 990 11155 1030 11195
rect 990 11075 1030 11115
rect 990 10995 1030 11035
rect 990 10915 1030 10955
rect 990 10835 1030 10875
rect 990 10755 1030 10795
rect 990 10675 1030 10715
rect 990 10595 1030 10635
rect 990 10515 1030 10555
rect 990 10435 1030 10475
rect 990 10355 1030 10395
rect 990 10275 1030 10315
rect 1105 12195 1145 12235
rect 1105 12115 1145 12155
rect 1105 12035 1145 12075
rect 1105 11955 1145 11995
rect 1105 11875 1145 11915
rect 1105 11795 1145 11835
rect 1105 11715 1145 11755
rect 1105 11635 1145 11675
rect 1105 11555 1145 11595
rect 1105 11475 1145 11515
rect 1105 11395 1145 11435
rect 1105 11315 1145 11355
rect 1105 11235 1145 11275
rect 1105 11155 1145 11195
rect 1105 11075 1145 11115
rect 1105 10995 1145 11035
rect 1105 10915 1145 10955
rect 1105 10835 1145 10875
rect 1105 10755 1145 10795
rect 1105 10675 1145 10715
rect 1105 10595 1145 10635
rect 1105 10515 1145 10555
rect 1105 10435 1145 10475
rect 1105 10355 1145 10395
rect 1105 10275 1145 10315
rect 1220 12195 1260 12235
rect 1220 12115 1260 12155
rect 1220 12035 1260 12075
rect 1220 11955 1260 11995
rect 1220 11875 1260 11915
rect 1220 11795 1260 11835
rect 1220 11715 1260 11755
rect 1220 11635 1260 11675
rect 1220 11555 1260 11595
rect 1220 11475 1260 11515
rect 1220 11395 1260 11435
rect 1220 11315 1260 11355
rect 1220 11235 1260 11275
rect 1220 11155 1260 11195
rect 1220 11075 1260 11115
rect 1220 10995 1260 11035
rect 1220 10915 1260 10955
rect 1220 10835 1260 10875
rect 1220 10755 1260 10795
rect 1220 10675 1260 10715
rect 1220 10595 1260 10635
rect 1220 10515 1260 10555
rect 1220 10435 1260 10475
rect 1220 10355 1260 10395
rect 1220 10275 1260 10315
rect 1335 12195 1375 12235
rect 1335 12115 1375 12155
rect 1335 12035 1375 12075
rect 1335 11955 1375 11995
rect 1335 11875 1375 11915
rect 1335 11795 1375 11835
rect 1335 11715 1375 11755
rect 1335 11635 1375 11675
rect 1335 11555 1375 11595
rect 1335 11475 1375 11515
rect 1335 11395 1375 11435
rect 1335 11315 1375 11355
rect 1335 11235 1375 11275
rect 1335 11155 1375 11195
rect 1335 11075 1375 11115
rect 1335 10995 1375 11035
rect 1335 10915 1375 10955
rect 1335 10835 1375 10875
rect 1335 10755 1375 10795
rect 1335 10675 1375 10715
rect 1335 10595 1375 10635
rect 1335 10515 1375 10555
rect 1335 10435 1375 10475
rect 1335 10355 1375 10395
rect 1335 10275 1375 10315
rect 1450 12195 1490 12235
rect 1450 12115 1490 12155
rect 1450 12035 1490 12075
rect 1450 11955 1490 11995
rect 1450 11875 1490 11915
rect 1450 11795 1490 11835
rect 1450 11715 1490 11755
rect 1450 11635 1490 11675
rect 1450 11555 1490 11595
rect 1450 11475 1490 11515
rect 1450 11395 1490 11435
rect 1450 11315 1490 11355
rect 1450 11235 1490 11275
rect 1450 11155 1490 11195
rect 1450 11075 1490 11115
rect 1450 10995 1490 11035
rect 1450 10915 1490 10955
rect 1450 10835 1490 10875
rect 1450 10755 1490 10795
rect 1450 10675 1490 10715
rect 1450 10595 1490 10635
rect 1450 10515 1490 10555
rect 1450 10435 1490 10475
rect 1450 10355 1490 10395
rect 1450 10275 1490 10315
rect 1565 12195 1605 12235
rect 1565 12115 1605 12155
rect 1565 12035 1605 12075
rect 1565 11955 1605 11995
rect 1565 11875 1605 11915
rect 1565 11795 1605 11835
rect 1565 11715 1605 11755
rect 1565 11635 1605 11675
rect 1565 11555 1605 11595
rect 1565 11475 1605 11515
rect 1565 11395 1605 11435
rect 1565 11315 1605 11355
rect 1565 11235 1605 11275
rect 1565 11155 1605 11195
rect 1565 11075 1605 11115
rect 1565 10995 1605 11035
rect 1565 10915 1605 10955
rect 1565 10835 1605 10875
rect 1565 10755 1605 10795
rect 1565 10675 1605 10715
rect 1565 10595 1605 10635
rect 1565 10515 1605 10555
rect 1565 10435 1605 10475
rect 1565 10355 1605 10395
rect 1565 10275 1605 10315
rect 1680 12195 1720 12235
rect 1680 12115 1720 12155
rect 1680 12035 1720 12075
rect 1680 11955 1720 11995
rect 1680 11875 1720 11915
rect 1680 11795 1720 11835
rect 1680 11715 1720 11755
rect 1680 11635 1720 11675
rect 1680 11555 1720 11595
rect 1680 11475 1720 11515
rect 1680 11395 1720 11435
rect 1680 11315 1720 11355
rect 1680 11235 1720 11275
rect 1680 11155 1720 11195
rect 1680 11075 1720 11115
rect 1680 10995 1720 11035
rect 1680 10915 1720 10955
rect 1680 10835 1720 10875
rect 1680 10755 1720 10795
rect 1680 10675 1720 10715
rect 1680 10595 1720 10635
rect 1680 10515 1720 10555
rect 1680 10435 1720 10475
rect 1680 10355 1720 10395
rect 1680 10275 1720 10315
rect 1795 12195 1835 12235
rect 1795 12115 1835 12155
rect 1795 12035 1835 12075
rect 1795 11955 1835 11995
rect 1795 11875 1835 11915
rect 1795 11795 1835 11835
rect 1795 11715 1835 11755
rect 1795 11635 1835 11675
rect 1795 11555 1835 11595
rect 1795 11475 1835 11515
rect 1795 11395 1835 11435
rect 1795 11315 1835 11355
rect 1795 11235 1835 11275
rect 1795 11155 1835 11195
rect 1795 11075 1835 11115
rect 1795 10995 1835 11035
rect 1795 10915 1835 10955
rect 1795 10835 1835 10875
rect 1795 10755 1835 10795
rect 1795 10675 1835 10715
rect 1795 10595 1835 10635
rect 1795 10515 1835 10555
rect 1795 10435 1835 10475
rect 1795 10355 1835 10395
rect 1795 10275 1835 10315
rect 1910 12195 1950 12235
rect 1910 12115 1950 12155
rect 1910 12035 1950 12075
rect 1910 11955 1950 11995
rect 1910 11875 1950 11915
rect 1910 11795 1950 11835
rect 1910 11715 1950 11755
rect 1910 11635 1950 11675
rect 1910 11555 1950 11595
rect 1910 11475 1950 11515
rect 1910 11395 1950 11435
rect 1910 11315 1950 11355
rect 1910 11235 1950 11275
rect 1910 11155 1950 11195
rect 1910 11075 1950 11115
rect 1910 10995 1950 11035
rect 1910 10915 1950 10955
rect 1910 10835 1950 10875
rect 1910 10755 1950 10795
rect 1910 10675 1950 10715
rect 1910 10595 1950 10635
rect 1910 10515 1950 10555
rect 1910 10435 1950 10475
rect 1910 10355 1950 10395
rect 1910 10275 1950 10315
rect 2025 12195 2065 12235
rect 2025 12115 2065 12155
rect 2025 12035 2065 12075
rect 2025 11955 2065 11995
rect 2025 11875 2065 11915
rect 2025 11795 2065 11835
rect 2025 11715 2065 11755
rect 2025 11635 2065 11675
rect 2025 11555 2065 11595
rect 2025 11475 2065 11515
rect 2025 11395 2065 11435
rect 2025 11315 2065 11355
rect 2025 11235 2065 11275
rect 2025 11155 2065 11195
rect 2025 11075 2065 11115
rect 2025 10995 2065 11035
rect 2025 10915 2065 10955
rect 2025 10835 2065 10875
rect 2025 10755 2065 10795
rect 2025 10675 2065 10715
rect 2025 10595 2065 10635
rect 2025 10515 2065 10555
rect 2025 10435 2065 10475
rect 2025 10355 2065 10395
rect 2025 10275 2065 10315
rect 2140 12195 2180 12235
rect 2140 12115 2180 12155
rect 2140 12035 2180 12075
rect 2140 11955 2180 11995
rect 2140 11875 2180 11915
rect 2140 11795 2180 11835
rect 2140 11715 2180 11755
rect 2140 11635 2180 11675
rect 2140 11555 2180 11595
rect 2140 11475 2180 11515
rect 2140 11395 2180 11435
rect 2140 11315 2180 11355
rect 2140 11235 2180 11275
rect 2140 11155 2180 11195
rect 2140 11075 2180 11115
rect 2140 10995 2180 11035
rect 2140 10915 2180 10955
rect 2140 10835 2180 10875
rect 2140 10755 2180 10795
rect 2140 10675 2180 10715
rect 2140 10595 2180 10635
rect 2140 10515 2180 10555
rect 2140 10435 2180 10475
rect 2140 10355 2180 10395
rect 2140 10275 2180 10315
rect 2255 12195 2295 12235
rect 2255 12115 2295 12155
rect 2255 12035 2295 12075
rect 2255 11955 2295 11995
rect 2255 11875 2295 11915
rect 2255 11795 2295 11835
rect 2255 11715 2295 11755
rect 2255 11635 2295 11675
rect 2255 11555 2295 11595
rect 2255 11475 2295 11515
rect 2255 11395 2295 11435
rect 2255 11315 2295 11355
rect 2255 11235 2295 11275
rect 2255 11155 2295 11195
rect 2255 11075 2295 11115
rect 2255 10995 2295 11035
rect 2255 10915 2295 10955
rect 2255 10835 2295 10875
rect 2255 10755 2295 10795
rect 2255 10675 2295 10715
rect 2255 10595 2295 10635
rect 2255 10515 2295 10555
rect 2255 10435 2295 10475
rect 2255 10355 2295 10395
rect 2255 10275 2295 10315
rect 2370 12195 2410 12235
rect 2370 12115 2410 12155
rect 2370 12035 2410 12075
rect 2370 11955 2410 11995
rect 2370 11875 2410 11915
rect 2370 11795 2410 11835
rect 2370 11715 2410 11755
rect 2370 11635 2410 11675
rect 2370 11555 2410 11595
rect 2370 11475 2410 11515
rect 2370 11395 2410 11435
rect 2370 11315 2410 11355
rect 2370 11235 2410 11275
rect 2370 11155 2410 11195
rect 2370 11075 2410 11115
rect 2370 10995 2410 11035
rect 2370 10915 2410 10955
rect 2370 10835 2410 10875
rect 2370 10755 2410 10795
rect 2370 10675 2410 10715
rect 2370 10595 2410 10635
rect 2370 10515 2410 10555
rect 2370 10435 2410 10475
rect 2370 10355 2410 10395
rect 2370 10275 2410 10315
rect 2485 12195 2525 12235
rect 2485 12115 2525 12155
rect 2485 12035 2525 12075
rect 2485 11955 2525 11995
rect 2485 11875 2525 11915
rect 2485 11795 2525 11835
rect 2485 11715 2525 11755
rect 2485 11635 2525 11675
rect 2485 11555 2525 11595
rect 2485 11475 2525 11515
rect 2485 11395 2525 11435
rect 2485 11315 2525 11355
rect 2485 11235 2525 11275
rect 2485 11155 2525 11195
rect 2485 11075 2525 11115
rect 2485 10995 2525 11035
rect 2485 10915 2525 10955
rect 2485 10835 2525 10875
rect 2485 10755 2525 10795
rect 2485 10675 2525 10715
rect 2485 10595 2525 10635
rect 2485 10515 2525 10555
rect 2485 10435 2525 10475
rect 2485 10355 2525 10395
rect 2485 10275 2525 10315
<< nsubdiff >>
rect -620 12475 880 12505
rect -620 12435 -390 12475
rect -350 12435 -230 12475
rect -190 12435 -70 12475
rect -30 12435 90 12475
rect 130 12435 250 12475
rect 290 12435 410 12475
rect 450 12435 570 12475
rect 610 12435 730 12475
rect 770 12435 880 12475
rect -620 12405 880 12435
rect 1265 12475 2755 12505
rect 1265 12435 1290 12475
rect 1330 12435 1450 12475
rect 1490 12435 1610 12475
rect 1650 12435 1770 12475
rect 1810 12435 1930 12475
rect 1970 12435 2090 12475
rect 2130 12435 2250 12475
rect 2290 12435 2410 12475
rect 2450 12435 2755 12475
rect -620 12235 -520 12405
rect 1265 12405 2755 12435
rect -620 12195 -590 12235
rect -550 12195 -520 12235
rect -620 12075 -520 12195
rect -620 12035 -590 12075
rect -550 12035 -520 12075
rect -620 11915 -520 12035
rect -620 11875 -590 11915
rect -550 11875 -520 11915
rect -620 11755 -520 11875
rect -620 11715 -590 11755
rect -550 11715 -520 11755
rect -620 11595 -520 11715
rect -620 11555 -590 11595
rect -550 11555 -520 11595
rect -620 11435 -520 11555
rect -620 11395 -590 11435
rect -550 11395 -520 11435
rect -620 11275 -520 11395
rect -620 11235 -590 11275
rect -550 11235 -520 11275
rect -620 11115 -520 11235
rect -620 11075 -590 11115
rect -550 11075 -520 11115
rect -620 10955 -520 11075
rect -620 10915 -590 10955
rect -550 10915 -520 10955
rect -620 10795 -520 10915
rect -620 10755 -590 10795
rect -550 10755 -520 10795
rect -620 10635 -520 10755
rect -620 10595 -590 10635
rect -550 10595 -520 10635
rect -620 10475 -520 10595
rect -620 10435 -590 10475
rect -550 10435 -520 10475
rect -620 10315 -520 10435
rect -620 10275 -590 10315
rect -550 10275 -520 10315
rect -620 10060 -520 10275
rect 2655 12155 2755 12405
rect 2655 12115 2685 12155
rect 2725 12115 2755 12155
rect 2655 11995 2755 12115
rect 2655 11955 2685 11995
rect 2725 11955 2755 11995
rect 2655 11835 2755 11955
rect 2655 11795 2685 11835
rect 2725 11795 2755 11835
rect 2655 11675 2755 11795
rect 2655 11635 2685 11675
rect 2725 11635 2755 11675
rect 2655 11515 2755 11635
rect 2655 11475 2685 11515
rect 2725 11475 2755 11515
rect 2655 11355 2755 11475
rect 2655 11315 2685 11355
rect 2725 11315 2755 11355
rect 2655 11195 2755 11315
rect 2655 11155 2685 11195
rect 2725 11155 2755 11195
rect 2655 10955 2755 11155
rect 2655 10915 2685 10955
rect 2725 10915 2755 10955
rect 2655 10795 2755 10915
rect 2655 10755 2685 10795
rect 2725 10755 2755 10795
rect 2655 10635 2755 10755
rect 2655 10595 2685 10635
rect 2725 10595 2755 10635
rect 2655 10475 2755 10595
rect 2655 10435 2685 10475
rect 2725 10435 2755 10475
rect 2655 10315 2755 10435
rect 2655 10275 2685 10315
rect 2725 10275 2755 10315
rect -620 10030 880 10060
rect 2655 10060 2755 10275
rect -620 9990 -390 10030
rect -350 9990 -230 10030
rect -190 9990 -70 10030
rect -30 9990 90 10030
rect 130 9990 250 10030
rect 290 9990 410 10030
rect 450 9990 570 10030
rect 610 9990 730 10030
rect 770 9990 880 10030
rect -620 9960 880 9990
rect 1260 10030 2755 10060
rect 1260 9990 1290 10030
rect 1330 9990 1450 10030
rect 1490 9990 1610 10030
rect 1650 9990 1770 10030
rect 1810 9990 1930 10030
rect 1970 9990 2090 10030
rect 2130 9990 2250 10030
rect 2290 9990 2410 10030
rect 2450 9990 2755 10030
rect 1260 9960 2755 9990
<< nsubdiffcont >>
rect -390 12435 -350 12475
rect -230 12435 -190 12475
rect -70 12435 -30 12475
rect 90 12435 130 12475
rect 250 12435 290 12475
rect 410 12435 450 12475
rect 570 12435 610 12475
rect 730 12435 770 12475
rect 1290 12435 1330 12475
rect 1450 12435 1490 12475
rect 1610 12435 1650 12475
rect 1770 12435 1810 12475
rect 1930 12435 1970 12475
rect 2090 12435 2130 12475
rect 2250 12435 2290 12475
rect 2410 12435 2450 12475
rect -590 12195 -550 12235
rect -590 12035 -550 12075
rect -590 11875 -550 11915
rect -590 11715 -550 11755
rect -590 11555 -550 11595
rect -590 11395 -550 11435
rect -590 11235 -550 11275
rect -590 11075 -550 11115
rect -590 10915 -550 10955
rect -590 10755 -550 10795
rect -590 10595 -550 10635
rect -590 10435 -550 10475
rect -590 10275 -550 10315
rect 2685 12115 2725 12155
rect 2685 11955 2725 11995
rect 2685 11795 2725 11835
rect 2685 11635 2725 11675
rect 2685 11475 2725 11515
rect 2685 11315 2725 11355
rect 2685 11155 2725 11195
rect 2685 10915 2725 10955
rect 2685 10755 2725 10795
rect 2685 10595 2725 10635
rect 2685 10435 2725 10475
rect 2685 10275 2725 10315
rect -390 9990 -350 10030
rect -230 9990 -190 10030
rect -70 9990 -30 10030
rect 90 9990 130 10030
rect 250 9990 290 10030
rect 410 9990 450 10030
rect 570 9990 610 10030
rect 730 9990 770 10030
rect 1290 9990 1330 10030
rect 1450 9990 1490 10030
rect 1610 9990 1650 10030
rect 1770 9990 1810 10030
rect 1930 9990 1970 10030
rect 2090 9990 2130 10030
rect 2250 9990 2290 10030
rect 2410 9990 2450 10030
<< poly >>
rect 1025 12490 1110 12505
rect 1025 12440 1040 12490
rect 1095 12440 1110 12490
rect 1025 12425 1110 12440
rect 1060 12320 1075 12425
rect -320 12305 2455 12320
rect -320 12270 -305 12305
rect -205 12270 -190 12305
rect -90 12270 -75 12305
rect 25 12270 40 12305
rect 140 12270 155 12305
rect 255 12270 270 12305
rect 370 12270 385 12305
rect 485 12270 500 12305
rect 600 12270 615 12305
rect 715 12270 730 12305
rect 830 12270 845 12305
rect 945 12270 960 12305
rect 1060 12270 1075 12305
rect 1175 12270 1190 12305
rect 1290 12270 1305 12305
rect 1405 12270 1420 12305
rect 1520 12270 1535 12305
rect 1635 12270 1650 12305
rect 1750 12270 1765 12305
rect 1865 12270 1880 12305
rect 1980 12270 1995 12305
rect 2095 12270 2110 12305
rect 2210 12270 2225 12305
rect 2325 12270 2340 12305
rect 2440 12270 2455 12305
rect -320 10200 -305 10245
rect -205 10200 -190 10245
rect -90 10200 -75 10245
rect 25 10200 40 10245
rect 140 10200 155 10245
rect 255 10200 270 10245
rect 370 10200 385 10245
rect 485 10200 500 10245
rect 600 10200 615 10245
rect 715 10200 730 10245
rect 830 10200 845 10245
rect 945 10200 960 10245
rect 1060 10200 1075 10245
rect 1175 10200 1190 10245
rect 1290 10200 1305 10245
rect 1405 10200 1420 10245
rect 1520 10200 1535 10245
rect 1635 10200 1650 10245
rect 1750 10200 1765 10245
rect 1865 10200 1880 10245
rect 1980 10200 1995 10245
rect 2095 10200 2110 10245
rect 2210 10200 2225 10245
rect 2325 10200 2340 10245
rect 2440 10200 2455 10245
rect -320 10185 2455 10200
rect 1060 10040 1075 10185
rect 1025 10025 1110 10040
rect 1025 9975 1040 10025
rect 1095 9975 1110 10025
rect 1025 9960 1110 9975
<< polycont >>
rect 1040 12440 1095 12490
rect 1040 9975 1095 10025
<< locali >>
rect 1025 12490 1110 12505
rect -405 12475 870 12490
rect -405 12435 -390 12475
rect -350 12435 -230 12475
rect -190 12435 -70 12475
rect -30 12435 90 12475
rect 130 12435 250 12475
rect 290 12435 410 12475
rect 450 12435 570 12475
rect 610 12435 730 12475
rect 770 12435 870 12475
rect -405 12420 870 12435
rect 1025 12440 1040 12490
rect 1095 12440 1110 12490
rect 1025 12425 1110 12440
rect 1275 12475 2545 12490
rect 1275 12435 1290 12475
rect 1330 12435 1450 12475
rect 1490 12435 1610 12475
rect 1650 12435 1770 12475
rect 1810 12435 1930 12475
rect 1970 12435 2090 12475
rect 2130 12435 2250 12475
rect 2290 12435 2410 12475
rect 2450 12435 2545 12475
rect 1275 12420 2545 12435
rect -605 12235 -535 12270
rect -605 12195 -590 12235
rect -550 12195 -535 12235
rect -605 12075 -535 12195
rect -605 12035 -590 12075
rect -550 12035 -535 12075
rect -605 11915 -535 12035
rect -605 11875 -590 11915
rect -550 11875 -535 11915
rect -605 11755 -535 11875
rect -605 11715 -590 11755
rect -550 11715 -535 11755
rect -605 11595 -535 11715
rect -605 11555 -590 11595
rect -550 11555 -535 11595
rect -605 11435 -535 11555
rect -605 11395 -590 11435
rect -550 11395 -535 11435
rect -605 11275 -535 11395
rect -605 11235 -590 11275
rect -550 11235 -535 11275
rect -605 11115 -535 11235
rect -605 11075 -590 11115
rect -550 11075 -535 11115
rect -605 10955 -535 11075
rect -605 10915 -590 10955
rect -550 10915 -535 10955
rect -605 10795 -535 10915
rect -605 10755 -590 10795
rect -550 10755 -535 10795
rect -605 10635 -535 10755
rect -605 10595 -590 10635
rect -550 10595 -535 10635
rect -605 10475 -535 10595
rect -605 10435 -590 10475
rect -550 10435 -535 10475
rect -605 10315 -535 10435
rect -605 10275 -590 10315
rect -550 10275 -535 10315
rect -605 10245 -535 10275
rect -405 12235 -334 12255
rect -405 12195 -390 12235
rect -350 12195 -334 12235
rect -405 12155 -334 12195
rect -405 12115 -390 12155
rect -350 12115 -334 12155
rect -405 12075 -334 12115
rect -405 12035 -390 12075
rect -350 12035 -334 12075
rect -405 11995 -334 12035
rect -405 11955 -390 11995
rect -350 11955 -334 11995
rect -405 11915 -334 11955
rect -405 11875 -390 11915
rect -350 11875 -334 11915
rect -405 11835 -334 11875
rect -405 11795 -390 11835
rect -350 11795 -334 11835
rect -405 11755 -334 11795
rect -405 11715 -390 11755
rect -350 11715 -334 11755
rect -405 11675 -334 11715
rect -405 11635 -390 11675
rect -350 11635 -334 11675
rect -405 11595 -334 11635
rect -405 11555 -390 11595
rect -350 11555 -334 11595
rect -405 11515 -334 11555
rect -405 11475 -390 11515
rect -350 11475 -334 11515
rect -405 11435 -334 11475
rect -405 11395 -390 11435
rect -350 11395 -334 11435
rect -405 11355 -334 11395
rect -405 11315 -390 11355
rect -350 11315 -334 11355
rect -405 11275 -334 11315
rect -405 11235 -390 11275
rect -350 11235 -334 11275
rect -405 11195 -334 11235
rect -405 11155 -390 11195
rect -350 11155 -334 11195
rect -405 11115 -334 11155
rect -405 11075 -390 11115
rect -350 11075 -334 11115
rect -405 11035 -334 11075
rect -405 10995 -390 11035
rect -350 10995 -334 11035
rect -405 10955 -334 10995
rect -405 10915 -390 10955
rect -350 10915 -334 10955
rect -405 10875 -334 10915
rect -405 10835 -390 10875
rect -350 10835 -334 10875
rect -405 10795 -334 10835
rect -405 10755 -390 10795
rect -350 10755 -334 10795
rect -405 10715 -334 10755
rect -405 10675 -390 10715
rect -350 10675 -334 10715
rect -405 10635 -334 10675
rect -405 10595 -390 10635
rect -350 10595 -334 10635
rect -405 10555 -334 10595
rect -405 10515 -390 10555
rect -350 10515 -334 10555
rect -405 10475 -334 10515
rect -405 10435 -390 10475
rect -350 10435 -334 10475
rect -405 10395 -334 10435
rect -405 10355 -390 10395
rect -350 10355 -334 10395
rect -405 10315 -334 10355
rect -405 10275 -390 10315
rect -350 10275 -334 10315
rect -405 10260 -334 10275
rect -290 12235 -220 12255
rect -290 12195 -275 12235
rect -235 12195 -220 12235
rect -290 12155 -220 12195
rect -290 12115 -275 12155
rect -235 12115 -220 12155
rect -290 12075 -220 12115
rect -290 12035 -275 12075
rect -235 12035 -220 12075
rect -290 11995 -220 12035
rect -290 11955 -275 11995
rect -235 11955 -220 11995
rect -290 11915 -220 11955
rect -290 11875 -275 11915
rect -235 11875 -220 11915
rect -290 11835 -220 11875
rect -290 11795 -275 11835
rect -235 11795 -220 11835
rect -290 11755 -220 11795
rect -290 11715 -275 11755
rect -235 11715 -220 11755
rect -290 11675 -220 11715
rect -290 11635 -275 11675
rect -235 11635 -220 11675
rect -290 11595 -220 11635
rect -290 11555 -275 11595
rect -235 11555 -220 11595
rect -290 11515 -220 11555
rect -290 11475 -275 11515
rect -235 11475 -220 11515
rect -290 11435 -220 11475
rect -290 11395 -275 11435
rect -235 11395 -220 11435
rect -290 11355 -220 11395
rect -290 11315 -275 11355
rect -235 11315 -220 11355
rect -290 11275 -220 11315
rect -290 11235 -275 11275
rect -235 11235 -220 11275
rect -290 11195 -220 11235
rect -290 11155 -275 11195
rect -235 11155 -220 11195
rect -290 11115 -220 11155
rect -290 11075 -275 11115
rect -235 11075 -220 11115
rect -290 11035 -220 11075
rect -290 10995 -275 11035
rect -235 10995 -220 11035
rect -290 10955 -220 10995
rect -290 10915 -275 10955
rect -235 10915 -220 10955
rect -290 10875 -220 10915
rect -290 10835 -275 10875
rect -235 10835 -220 10875
rect -290 10795 -220 10835
rect -290 10755 -275 10795
rect -235 10755 -220 10795
rect -290 10715 -220 10755
rect -290 10675 -275 10715
rect -235 10675 -220 10715
rect -290 10635 -220 10675
rect -290 10595 -275 10635
rect -235 10595 -220 10635
rect -290 10555 -220 10595
rect -290 10515 -275 10555
rect -235 10515 -220 10555
rect -290 10475 -220 10515
rect -290 10435 -275 10475
rect -235 10435 -220 10475
rect -290 10395 -220 10435
rect -290 10355 -275 10395
rect -235 10355 -220 10395
rect -290 10315 -220 10355
rect -290 10275 -275 10315
rect -235 10275 -220 10315
rect -290 10260 -220 10275
rect -175 12235 -105 12255
rect -175 12195 -160 12235
rect -120 12195 -105 12235
rect -175 12155 -105 12195
rect -175 12115 -160 12155
rect -120 12115 -105 12155
rect -175 12075 -105 12115
rect -175 12035 -160 12075
rect -120 12035 -105 12075
rect -175 11995 -105 12035
rect -175 11955 -160 11995
rect -120 11955 -105 11995
rect -175 11915 -105 11955
rect -175 11875 -160 11915
rect -120 11875 -105 11915
rect -175 11835 -105 11875
rect -175 11795 -160 11835
rect -120 11795 -105 11835
rect -175 11755 -105 11795
rect -175 11715 -160 11755
rect -120 11715 -105 11755
rect -175 11675 -105 11715
rect -175 11635 -160 11675
rect -120 11635 -105 11675
rect -175 11595 -105 11635
rect -175 11555 -160 11595
rect -120 11555 -105 11595
rect -175 11515 -105 11555
rect -175 11475 -160 11515
rect -120 11475 -105 11515
rect -175 11435 -105 11475
rect -175 11395 -160 11435
rect -120 11395 -105 11435
rect -175 11355 -105 11395
rect -175 11315 -160 11355
rect -120 11315 -105 11355
rect -175 11275 -105 11315
rect -175 11235 -160 11275
rect -120 11235 -105 11275
rect -175 11195 -105 11235
rect -175 11155 -160 11195
rect -120 11155 -105 11195
rect -175 11115 -105 11155
rect -175 11075 -160 11115
rect -120 11075 -105 11115
rect -175 11035 -105 11075
rect -175 10995 -160 11035
rect -120 10995 -105 11035
rect -175 10955 -105 10995
rect -175 10915 -160 10955
rect -120 10915 -105 10955
rect -175 10875 -105 10915
rect -175 10835 -160 10875
rect -120 10835 -105 10875
rect -175 10795 -105 10835
rect -175 10755 -160 10795
rect -120 10755 -105 10795
rect -175 10715 -105 10755
rect -175 10675 -160 10715
rect -120 10675 -105 10715
rect -175 10635 -105 10675
rect -175 10595 -160 10635
rect -120 10595 -105 10635
rect -175 10555 -105 10595
rect -175 10515 -160 10555
rect -120 10515 -105 10555
rect -175 10475 -105 10515
rect -175 10435 -160 10475
rect -120 10435 -105 10475
rect -175 10395 -105 10435
rect -175 10355 -160 10395
rect -120 10355 -105 10395
rect -175 10315 -105 10355
rect -175 10275 -160 10315
rect -120 10275 -105 10315
rect -175 10260 -105 10275
rect -60 12235 10 12255
rect -60 12195 -45 12235
rect -5 12195 10 12235
rect -60 12155 10 12195
rect -60 12115 -45 12155
rect -5 12115 10 12155
rect -60 12075 10 12115
rect -60 12035 -45 12075
rect -5 12035 10 12075
rect -60 11995 10 12035
rect -60 11955 -45 11995
rect -5 11955 10 11995
rect -60 11915 10 11955
rect -60 11875 -45 11915
rect -5 11875 10 11915
rect -60 11835 10 11875
rect -60 11795 -45 11835
rect -5 11795 10 11835
rect -60 11755 10 11795
rect -60 11715 -45 11755
rect -5 11715 10 11755
rect -60 11675 10 11715
rect -60 11635 -45 11675
rect -5 11635 10 11675
rect -60 11595 10 11635
rect -60 11555 -45 11595
rect -5 11555 10 11595
rect -60 11515 10 11555
rect -60 11475 -45 11515
rect -5 11475 10 11515
rect -60 11435 10 11475
rect -60 11395 -45 11435
rect -5 11395 10 11435
rect -60 11355 10 11395
rect -60 11315 -45 11355
rect -5 11315 10 11355
rect -60 11275 10 11315
rect -60 11235 -45 11275
rect -5 11235 10 11275
rect -60 11195 10 11235
rect -60 11155 -45 11195
rect -5 11155 10 11195
rect -60 11115 10 11155
rect -60 11075 -45 11115
rect -5 11075 10 11115
rect -60 11035 10 11075
rect -60 10995 -45 11035
rect -5 10995 10 11035
rect -60 10955 10 10995
rect -60 10915 -45 10955
rect -5 10915 10 10955
rect -60 10875 10 10915
rect -60 10835 -45 10875
rect -5 10835 10 10875
rect -60 10795 10 10835
rect -60 10755 -45 10795
rect -5 10755 10 10795
rect -60 10715 10 10755
rect -60 10675 -45 10715
rect -5 10675 10 10715
rect -60 10635 10 10675
rect -60 10595 -45 10635
rect -5 10595 10 10635
rect -60 10555 10 10595
rect -60 10515 -45 10555
rect -5 10515 10 10555
rect -60 10475 10 10515
rect -60 10435 -45 10475
rect -5 10435 10 10475
rect -60 10395 10 10435
rect -60 10355 -45 10395
rect -5 10355 10 10395
rect -60 10315 10 10355
rect -60 10275 -45 10315
rect -5 10275 10 10315
rect -60 10260 10 10275
rect 55 12235 125 12255
rect 55 12195 70 12235
rect 110 12195 125 12235
rect 55 12155 125 12195
rect 55 12115 70 12155
rect 110 12115 125 12155
rect 55 12075 125 12115
rect 55 12035 70 12075
rect 110 12035 125 12075
rect 55 11995 125 12035
rect 55 11955 70 11995
rect 110 11955 125 11995
rect 55 11915 125 11955
rect 55 11875 70 11915
rect 110 11875 125 11915
rect 55 11835 125 11875
rect 55 11795 70 11835
rect 110 11795 125 11835
rect 55 11755 125 11795
rect 55 11715 70 11755
rect 110 11715 125 11755
rect 55 11675 125 11715
rect 55 11635 70 11675
rect 110 11635 125 11675
rect 55 11595 125 11635
rect 55 11555 70 11595
rect 110 11555 125 11595
rect 55 11515 125 11555
rect 55 11475 70 11515
rect 110 11475 125 11515
rect 55 11435 125 11475
rect 55 11395 70 11435
rect 110 11395 125 11435
rect 55 11355 125 11395
rect 55 11315 70 11355
rect 110 11315 125 11355
rect 55 11275 125 11315
rect 55 11235 70 11275
rect 110 11235 125 11275
rect 55 11195 125 11235
rect 55 11155 70 11195
rect 110 11155 125 11195
rect 55 11115 125 11155
rect 55 11075 70 11115
rect 110 11075 125 11115
rect 55 11035 125 11075
rect 55 10995 70 11035
rect 110 10995 125 11035
rect 55 10955 125 10995
rect 55 10915 70 10955
rect 110 10915 125 10955
rect 55 10875 125 10915
rect 55 10835 70 10875
rect 110 10835 125 10875
rect 55 10795 125 10835
rect 55 10755 70 10795
rect 110 10755 125 10795
rect 55 10715 125 10755
rect 55 10675 70 10715
rect 110 10675 125 10715
rect 55 10635 125 10675
rect 55 10595 70 10635
rect 110 10595 125 10635
rect 55 10555 125 10595
rect 55 10515 70 10555
rect 110 10515 125 10555
rect 55 10475 125 10515
rect 55 10435 70 10475
rect 110 10435 125 10475
rect 55 10395 125 10435
rect 55 10355 70 10395
rect 110 10355 125 10395
rect 55 10315 125 10355
rect 55 10275 70 10315
rect 110 10275 125 10315
rect 55 10260 125 10275
rect 170 12235 240 12255
rect 170 12195 185 12235
rect 225 12195 240 12235
rect 170 12155 240 12195
rect 170 12115 185 12155
rect 225 12115 240 12155
rect 170 12075 240 12115
rect 170 12035 185 12075
rect 225 12035 240 12075
rect 170 11995 240 12035
rect 170 11955 185 11995
rect 225 11955 240 11995
rect 170 11915 240 11955
rect 170 11875 185 11915
rect 225 11875 240 11915
rect 170 11835 240 11875
rect 170 11795 185 11835
rect 225 11795 240 11835
rect 170 11755 240 11795
rect 170 11715 185 11755
rect 225 11715 240 11755
rect 170 11675 240 11715
rect 170 11635 185 11675
rect 225 11635 240 11675
rect 170 11595 240 11635
rect 170 11555 185 11595
rect 225 11555 240 11595
rect 170 11515 240 11555
rect 170 11475 185 11515
rect 225 11475 240 11515
rect 170 11435 240 11475
rect 170 11395 185 11435
rect 225 11395 240 11435
rect 170 11355 240 11395
rect 170 11315 185 11355
rect 225 11315 240 11355
rect 170 11275 240 11315
rect 170 11235 185 11275
rect 225 11235 240 11275
rect 170 11195 240 11235
rect 170 11155 185 11195
rect 225 11155 240 11195
rect 170 11115 240 11155
rect 170 11075 185 11115
rect 225 11075 240 11115
rect 170 11035 240 11075
rect 170 10995 185 11035
rect 225 10995 240 11035
rect 170 10955 240 10995
rect 170 10915 185 10955
rect 225 10915 240 10955
rect 170 10875 240 10915
rect 170 10835 185 10875
rect 225 10835 240 10875
rect 170 10795 240 10835
rect 170 10755 185 10795
rect 225 10755 240 10795
rect 170 10715 240 10755
rect 170 10675 185 10715
rect 225 10675 240 10715
rect 170 10635 240 10675
rect 170 10595 185 10635
rect 225 10595 240 10635
rect 170 10555 240 10595
rect 170 10515 185 10555
rect 225 10515 240 10555
rect 170 10475 240 10515
rect 170 10435 185 10475
rect 225 10435 240 10475
rect 170 10395 240 10435
rect 170 10355 185 10395
rect 225 10355 240 10395
rect 170 10315 240 10355
rect 170 10275 185 10315
rect 225 10275 240 10315
rect 170 10260 240 10275
rect 285 12235 355 12255
rect 285 12195 300 12235
rect 340 12195 355 12235
rect 285 12155 355 12195
rect 285 12115 300 12155
rect 340 12115 355 12155
rect 285 12075 355 12115
rect 285 12035 300 12075
rect 340 12035 355 12075
rect 285 11995 355 12035
rect 285 11955 300 11995
rect 340 11955 355 11995
rect 285 11915 355 11955
rect 285 11875 300 11915
rect 340 11875 355 11915
rect 285 11835 355 11875
rect 285 11795 300 11835
rect 340 11795 355 11835
rect 285 11755 355 11795
rect 285 11715 300 11755
rect 340 11715 355 11755
rect 285 11675 355 11715
rect 285 11635 300 11675
rect 340 11635 355 11675
rect 285 11595 355 11635
rect 285 11555 300 11595
rect 340 11555 355 11595
rect 285 11515 355 11555
rect 285 11475 300 11515
rect 340 11475 355 11515
rect 285 11435 355 11475
rect 285 11395 300 11435
rect 340 11395 355 11435
rect 285 11355 355 11395
rect 285 11315 300 11355
rect 340 11315 355 11355
rect 285 11275 355 11315
rect 285 11235 300 11275
rect 340 11235 355 11275
rect 285 11195 355 11235
rect 285 11155 300 11195
rect 340 11155 355 11195
rect 285 11115 355 11155
rect 285 11075 300 11115
rect 340 11075 355 11115
rect 285 11035 355 11075
rect 285 10995 300 11035
rect 340 10995 355 11035
rect 285 10955 355 10995
rect 285 10915 300 10955
rect 340 10915 355 10955
rect 285 10875 355 10915
rect 285 10835 300 10875
rect 340 10835 355 10875
rect 285 10795 355 10835
rect 285 10755 300 10795
rect 340 10755 355 10795
rect 285 10715 355 10755
rect 285 10675 300 10715
rect 340 10675 355 10715
rect 285 10635 355 10675
rect 285 10595 300 10635
rect 340 10595 355 10635
rect 285 10555 355 10595
rect 285 10515 300 10555
rect 340 10515 355 10555
rect 285 10475 355 10515
rect 285 10435 300 10475
rect 340 10435 355 10475
rect 285 10395 355 10435
rect 285 10355 300 10395
rect 340 10355 355 10395
rect 285 10315 355 10355
rect 285 10275 300 10315
rect 340 10275 355 10315
rect 285 10260 355 10275
rect 400 12235 470 12255
rect 400 12195 415 12235
rect 455 12195 470 12235
rect 400 12155 470 12195
rect 400 12115 415 12155
rect 455 12115 470 12155
rect 400 12075 470 12115
rect 400 12035 415 12075
rect 455 12035 470 12075
rect 400 11995 470 12035
rect 400 11955 415 11995
rect 455 11955 470 11995
rect 400 11915 470 11955
rect 400 11875 415 11915
rect 455 11875 470 11915
rect 400 11835 470 11875
rect 400 11795 415 11835
rect 455 11795 470 11835
rect 400 11755 470 11795
rect 400 11715 415 11755
rect 455 11715 470 11755
rect 400 11675 470 11715
rect 400 11635 415 11675
rect 455 11635 470 11675
rect 400 11595 470 11635
rect 400 11555 415 11595
rect 455 11555 470 11595
rect 400 11515 470 11555
rect 400 11475 415 11515
rect 455 11475 470 11515
rect 400 11435 470 11475
rect 400 11395 415 11435
rect 455 11395 470 11435
rect 400 11355 470 11395
rect 400 11315 415 11355
rect 455 11315 470 11355
rect 400 11275 470 11315
rect 400 11235 415 11275
rect 455 11235 470 11275
rect 400 11195 470 11235
rect 400 11155 415 11195
rect 455 11155 470 11195
rect 400 11115 470 11155
rect 400 11075 415 11115
rect 455 11075 470 11115
rect 400 11035 470 11075
rect 400 10995 415 11035
rect 455 10995 470 11035
rect 400 10955 470 10995
rect 400 10915 415 10955
rect 455 10915 470 10955
rect 400 10875 470 10915
rect 400 10835 415 10875
rect 455 10835 470 10875
rect 400 10795 470 10835
rect 400 10755 415 10795
rect 455 10755 470 10795
rect 400 10715 470 10755
rect 400 10675 415 10715
rect 455 10675 470 10715
rect 400 10635 470 10675
rect 400 10595 415 10635
rect 455 10595 470 10635
rect 400 10555 470 10595
rect 400 10515 415 10555
rect 455 10515 470 10555
rect 400 10475 470 10515
rect 400 10435 415 10475
rect 455 10435 470 10475
rect 400 10395 470 10435
rect 400 10355 415 10395
rect 455 10355 470 10395
rect 400 10315 470 10355
rect 400 10275 415 10315
rect 455 10275 470 10315
rect 400 10260 470 10275
rect 515 12235 585 12255
rect 515 12195 530 12235
rect 570 12195 585 12235
rect 515 12155 585 12195
rect 515 12115 530 12155
rect 570 12115 585 12155
rect 515 12075 585 12115
rect 515 12035 530 12075
rect 570 12035 585 12075
rect 515 11995 585 12035
rect 515 11955 530 11995
rect 570 11955 585 11995
rect 515 11915 585 11955
rect 515 11875 530 11915
rect 570 11875 585 11915
rect 515 11835 585 11875
rect 515 11795 530 11835
rect 570 11795 585 11835
rect 515 11755 585 11795
rect 515 11715 530 11755
rect 570 11715 585 11755
rect 515 11675 585 11715
rect 515 11635 530 11675
rect 570 11635 585 11675
rect 515 11595 585 11635
rect 515 11555 530 11595
rect 570 11555 585 11595
rect 515 11515 585 11555
rect 515 11475 530 11515
rect 570 11475 585 11515
rect 515 11435 585 11475
rect 515 11395 530 11435
rect 570 11395 585 11435
rect 515 11355 585 11395
rect 515 11315 530 11355
rect 570 11315 585 11355
rect 515 11275 585 11315
rect 515 11235 530 11275
rect 570 11235 585 11275
rect 515 11195 585 11235
rect 515 11155 530 11195
rect 570 11155 585 11195
rect 515 11115 585 11155
rect 515 11075 530 11115
rect 570 11075 585 11115
rect 515 11035 585 11075
rect 515 10995 530 11035
rect 570 10995 585 11035
rect 515 10955 585 10995
rect 515 10915 530 10955
rect 570 10915 585 10955
rect 515 10875 585 10915
rect 515 10835 530 10875
rect 570 10835 585 10875
rect 515 10795 585 10835
rect 515 10755 530 10795
rect 570 10755 585 10795
rect 515 10715 585 10755
rect 515 10675 530 10715
rect 570 10675 585 10715
rect 515 10635 585 10675
rect 515 10595 530 10635
rect 570 10595 585 10635
rect 515 10555 585 10595
rect 515 10515 530 10555
rect 570 10515 585 10555
rect 515 10475 585 10515
rect 515 10435 530 10475
rect 570 10435 585 10475
rect 515 10395 585 10435
rect 515 10355 530 10395
rect 570 10355 585 10395
rect 515 10315 585 10355
rect 515 10275 530 10315
rect 570 10275 585 10315
rect 515 10260 585 10275
rect 630 12235 700 12255
rect 630 12195 645 12235
rect 685 12195 700 12235
rect 630 12155 700 12195
rect 630 12115 645 12155
rect 685 12115 700 12155
rect 630 12075 700 12115
rect 630 12035 645 12075
rect 685 12035 700 12075
rect 630 11995 700 12035
rect 630 11955 645 11995
rect 685 11955 700 11995
rect 630 11915 700 11955
rect 630 11875 645 11915
rect 685 11875 700 11915
rect 630 11835 700 11875
rect 630 11795 645 11835
rect 685 11795 700 11835
rect 630 11755 700 11795
rect 630 11715 645 11755
rect 685 11715 700 11755
rect 630 11675 700 11715
rect 630 11635 645 11675
rect 685 11635 700 11675
rect 630 11595 700 11635
rect 630 11555 645 11595
rect 685 11555 700 11595
rect 630 11515 700 11555
rect 630 11475 645 11515
rect 685 11475 700 11515
rect 630 11435 700 11475
rect 630 11395 645 11435
rect 685 11395 700 11435
rect 630 11355 700 11395
rect 630 11315 645 11355
rect 685 11315 700 11355
rect 630 11275 700 11315
rect 630 11235 645 11275
rect 685 11235 700 11275
rect 630 11195 700 11235
rect 630 11155 645 11195
rect 685 11155 700 11195
rect 630 11115 700 11155
rect 630 11075 645 11115
rect 685 11075 700 11115
rect 630 11035 700 11075
rect 630 10995 645 11035
rect 685 10995 700 11035
rect 630 10955 700 10995
rect 630 10915 645 10955
rect 685 10915 700 10955
rect 630 10875 700 10915
rect 630 10835 645 10875
rect 685 10835 700 10875
rect 630 10795 700 10835
rect 630 10755 645 10795
rect 685 10755 700 10795
rect 630 10715 700 10755
rect 630 10675 645 10715
rect 685 10675 700 10715
rect 630 10635 700 10675
rect 630 10595 645 10635
rect 685 10595 700 10635
rect 630 10555 700 10595
rect 630 10515 645 10555
rect 685 10515 700 10555
rect 630 10475 700 10515
rect 630 10435 645 10475
rect 685 10435 700 10475
rect 630 10395 700 10435
rect 630 10355 645 10395
rect 685 10355 700 10395
rect 630 10315 700 10355
rect 630 10275 645 10315
rect 685 10275 700 10315
rect 630 10260 700 10275
rect 745 12235 815 12255
rect 745 12195 760 12235
rect 800 12195 815 12235
rect 745 12155 815 12195
rect 745 12115 760 12155
rect 800 12115 815 12155
rect 745 12075 815 12115
rect 745 12035 760 12075
rect 800 12035 815 12075
rect 745 11995 815 12035
rect 745 11955 760 11995
rect 800 11955 815 11995
rect 745 11915 815 11955
rect 745 11875 760 11915
rect 800 11875 815 11915
rect 745 11835 815 11875
rect 745 11795 760 11835
rect 800 11795 815 11835
rect 745 11755 815 11795
rect 745 11715 760 11755
rect 800 11715 815 11755
rect 745 11675 815 11715
rect 745 11635 760 11675
rect 800 11635 815 11675
rect 745 11595 815 11635
rect 745 11555 760 11595
rect 800 11555 815 11595
rect 745 11515 815 11555
rect 745 11475 760 11515
rect 800 11475 815 11515
rect 745 11435 815 11475
rect 745 11395 760 11435
rect 800 11395 815 11435
rect 745 11355 815 11395
rect 745 11315 760 11355
rect 800 11315 815 11355
rect 745 11275 815 11315
rect 745 11235 760 11275
rect 800 11235 815 11275
rect 745 11195 815 11235
rect 745 11155 760 11195
rect 800 11155 815 11195
rect 745 11115 815 11155
rect 745 11075 760 11115
rect 800 11075 815 11115
rect 745 11035 815 11075
rect 745 10995 760 11035
rect 800 10995 815 11035
rect 745 10955 815 10995
rect 745 10915 760 10955
rect 800 10915 815 10955
rect 745 10875 815 10915
rect 745 10835 760 10875
rect 800 10835 815 10875
rect 745 10795 815 10835
rect 745 10755 760 10795
rect 800 10755 815 10795
rect 745 10715 815 10755
rect 745 10675 760 10715
rect 800 10675 815 10715
rect 745 10635 815 10675
rect 745 10595 760 10635
rect 800 10595 815 10635
rect 745 10555 815 10595
rect 745 10515 760 10555
rect 800 10515 815 10555
rect 745 10475 815 10515
rect 745 10435 760 10475
rect 800 10435 815 10475
rect 745 10395 815 10435
rect 745 10355 760 10395
rect 800 10355 815 10395
rect 745 10315 815 10355
rect 745 10275 760 10315
rect 800 10275 815 10315
rect 745 10260 815 10275
rect 860 12235 930 12255
rect 860 12195 875 12235
rect 915 12195 930 12235
rect 860 12155 930 12195
rect 860 12115 875 12155
rect 915 12115 930 12155
rect 860 12075 930 12115
rect 860 12035 875 12075
rect 915 12035 930 12075
rect 860 11995 930 12035
rect 860 11955 875 11995
rect 915 11955 930 11995
rect 860 11915 930 11955
rect 860 11875 875 11915
rect 915 11875 930 11915
rect 860 11835 930 11875
rect 860 11795 875 11835
rect 915 11795 930 11835
rect 860 11755 930 11795
rect 860 11715 875 11755
rect 915 11715 930 11755
rect 860 11675 930 11715
rect 860 11635 875 11675
rect 915 11635 930 11675
rect 860 11595 930 11635
rect 860 11555 875 11595
rect 915 11555 930 11595
rect 860 11515 930 11555
rect 860 11475 875 11515
rect 915 11475 930 11515
rect 860 11435 930 11475
rect 860 11395 875 11435
rect 915 11395 930 11435
rect 860 11355 930 11395
rect 860 11315 875 11355
rect 915 11315 930 11355
rect 860 11275 930 11315
rect 860 11235 875 11275
rect 915 11235 930 11275
rect 860 11195 930 11235
rect 860 11155 875 11195
rect 915 11155 930 11195
rect 860 11115 930 11155
rect 860 11075 875 11115
rect 915 11075 930 11115
rect 860 11035 930 11075
rect 860 10995 875 11035
rect 915 10995 930 11035
rect 860 10955 930 10995
rect 860 10915 875 10955
rect 915 10915 930 10955
rect 860 10875 930 10915
rect 860 10835 875 10875
rect 915 10835 930 10875
rect 860 10795 930 10835
rect 860 10755 875 10795
rect 915 10755 930 10795
rect 860 10715 930 10755
rect 860 10675 875 10715
rect 915 10675 930 10715
rect 860 10635 930 10675
rect 860 10595 875 10635
rect 915 10595 930 10635
rect 860 10555 930 10595
rect 860 10515 875 10555
rect 915 10515 930 10555
rect 860 10475 930 10515
rect 860 10435 875 10475
rect 915 10435 930 10475
rect 860 10395 930 10435
rect 860 10355 875 10395
rect 915 10355 930 10395
rect 860 10315 930 10355
rect 860 10275 875 10315
rect 915 10275 930 10315
rect 860 10260 930 10275
rect 975 12235 1045 12255
rect 975 12195 990 12235
rect 1030 12195 1045 12235
rect 975 12155 1045 12195
rect 975 12115 990 12155
rect 1030 12115 1045 12155
rect 975 12075 1045 12115
rect 975 12035 990 12075
rect 1030 12035 1045 12075
rect 975 11995 1045 12035
rect 975 11955 990 11995
rect 1030 11955 1045 11995
rect 975 11915 1045 11955
rect 975 11875 990 11915
rect 1030 11875 1045 11915
rect 975 11835 1045 11875
rect 975 11795 990 11835
rect 1030 11795 1045 11835
rect 975 11755 1045 11795
rect 975 11715 990 11755
rect 1030 11715 1045 11755
rect 975 11675 1045 11715
rect 975 11635 990 11675
rect 1030 11635 1045 11675
rect 975 11595 1045 11635
rect 975 11555 990 11595
rect 1030 11555 1045 11595
rect 975 11515 1045 11555
rect 975 11475 990 11515
rect 1030 11475 1045 11515
rect 975 11435 1045 11475
rect 975 11395 990 11435
rect 1030 11395 1045 11435
rect 975 11355 1045 11395
rect 975 11315 990 11355
rect 1030 11315 1045 11355
rect 975 11275 1045 11315
rect 975 11235 990 11275
rect 1030 11235 1045 11275
rect 975 11195 1045 11235
rect 975 11155 990 11195
rect 1030 11155 1045 11195
rect 975 11115 1045 11155
rect 975 11075 990 11115
rect 1030 11075 1045 11115
rect 975 11035 1045 11075
rect 975 10995 990 11035
rect 1030 10995 1045 11035
rect 975 10955 1045 10995
rect 975 10915 990 10955
rect 1030 10915 1045 10955
rect 975 10875 1045 10915
rect 975 10835 990 10875
rect 1030 10835 1045 10875
rect 975 10795 1045 10835
rect 975 10755 990 10795
rect 1030 10755 1045 10795
rect 975 10715 1045 10755
rect 975 10675 990 10715
rect 1030 10675 1045 10715
rect 975 10635 1045 10675
rect 975 10595 990 10635
rect 1030 10595 1045 10635
rect 975 10555 1045 10595
rect 975 10515 990 10555
rect 1030 10515 1045 10555
rect 975 10475 1045 10515
rect 975 10435 990 10475
rect 1030 10435 1045 10475
rect 975 10395 1045 10435
rect 975 10355 990 10395
rect 1030 10355 1045 10395
rect 975 10315 1045 10355
rect 975 10275 990 10315
rect 1030 10275 1045 10315
rect 975 10260 1045 10275
rect 1090 12235 1160 12255
rect 1090 12195 1105 12235
rect 1145 12195 1160 12235
rect 1090 12155 1160 12195
rect 1090 12115 1105 12155
rect 1145 12115 1160 12155
rect 1090 12075 1160 12115
rect 1090 12035 1105 12075
rect 1145 12035 1160 12075
rect 1090 11995 1160 12035
rect 1090 11955 1105 11995
rect 1145 11955 1160 11995
rect 1090 11915 1160 11955
rect 1090 11875 1105 11915
rect 1145 11875 1160 11915
rect 1090 11835 1160 11875
rect 1090 11795 1105 11835
rect 1145 11795 1160 11835
rect 1090 11755 1160 11795
rect 1090 11715 1105 11755
rect 1145 11715 1160 11755
rect 1090 11675 1160 11715
rect 1090 11635 1105 11675
rect 1145 11635 1160 11675
rect 1090 11595 1160 11635
rect 1090 11555 1105 11595
rect 1145 11555 1160 11595
rect 1090 11515 1160 11555
rect 1090 11475 1105 11515
rect 1145 11475 1160 11515
rect 1090 11435 1160 11475
rect 1090 11395 1105 11435
rect 1145 11395 1160 11435
rect 1090 11355 1160 11395
rect 1090 11315 1105 11355
rect 1145 11315 1160 11355
rect 1090 11275 1160 11315
rect 1090 11235 1105 11275
rect 1145 11235 1160 11275
rect 1090 11195 1160 11235
rect 1090 11155 1105 11195
rect 1145 11155 1160 11195
rect 1090 11115 1160 11155
rect 1090 11075 1105 11115
rect 1145 11075 1160 11115
rect 1090 11035 1160 11075
rect 1090 10995 1105 11035
rect 1145 10995 1160 11035
rect 1090 10955 1160 10995
rect 1090 10915 1105 10955
rect 1145 10915 1160 10955
rect 1090 10875 1160 10915
rect 1090 10835 1105 10875
rect 1145 10835 1160 10875
rect 1090 10795 1160 10835
rect 1090 10755 1105 10795
rect 1145 10755 1160 10795
rect 1090 10715 1160 10755
rect 1090 10675 1105 10715
rect 1145 10675 1160 10715
rect 1090 10635 1160 10675
rect 1090 10595 1105 10635
rect 1145 10595 1160 10635
rect 1090 10555 1160 10595
rect 1090 10515 1105 10555
rect 1145 10515 1160 10555
rect 1090 10475 1160 10515
rect 1090 10435 1105 10475
rect 1145 10435 1160 10475
rect 1090 10395 1160 10435
rect 1090 10355 1105 10395
rect 1145 10355 1160 10395
rect 1090 10315 1160 10355
rect 1090 10275 1105 10315
rect 1145 10275 1160 10315
rect 1090 10260 1160 10275
rect 1205 12235 1275 12255
rect 1205 12195 1220 12235
rect 1260 12195 1275 12235
rect 1205 12155 1275 12195
rect 1205 12115 1220 12155
rect 1260 12115 1275 12155
rect 1205 12075 1275 12115
rect 1205 12035 1220 12075
rect 1260 12035 1275 12075
rect 1205 11995 1275 12035
rect 1205 11955 1220 11995
rect 1260 11955 1275 11995
rect 1205 11915 1275 11955
rect 1205 11875 1220 11915
rect 1260 11875 1275 11915
rect 1205 11835 1275 11875
rect 1205 11795 1220 11835
rect 1260 11795 1275 11835
rect 1205 11755 1275 11795
rect 1205 11715 1220 11755
rect 1260 11715 1275 11755
rect 1205 11675 1275 11715
rect 1205 11635 1220 11675
rect 1260 11635 1275 11675
rect 1205 11595 1275 11635
rect 1205 11555 1220 11595
rect 1260 11555 1275 11595
rect 1205 11515 1275 11555
rect 1205 11475 1220 11515
rect 1260 11475 1275 11515
rect 1205 11435 1275 11475
rect 1205 11395 1220 11435
rect 1260 11395 1275 11435
rect 1205 11355 1275 11395
rect 1205 11315 1220 11355
rect 1260 11315 1275 11355
rect 1205 11275 1275 11315
rect 1205 11235 1220 11275
rect 1260 11235 1275 11275
rect 1205 11195 1275 11235
rect 1205 11155 1220 11195
rect 1260 11155 1275 11195
rect 1205 11115 1275 11155
rect 1205 11075 1220 11115
rect 1260 11075 1275 11115
rect 1205 11035 1275 11075
rect 1205 10995 1220 11035
rect 1260 10995 1275 11035
rect 1205 10955 1275 10995
rect 1205 10915 1220 10955
rect 1260 10915 1275 10955
rect 1205 10875 1275 10915
rect 1205 10835 1220 10875
rect 1260 10835 1275 10875
rect 1205 10795 1275 10835
rect 1205 10755 1220 10795
rect 1260 10755 1275 10795
rect 1205 10715 1275 10755
rect 1205 10675 1220 10715
rect 1260 10675 1275 10715
rect 1205 10635 1275 10675
rect 1205 10595 1220 10635
rect 1260 10595 1275 10635
rect 1205 10555 1275 10595
rect 1205 10515 1220 10555
rect 1260 10515 1275 10555
rect 1205 10475 1275 10515
rect 1205 10435 1220 10475
rect 1260 10435 1275 10475
rect 1205 10395 1275 10435
rect 1205 10355 1220 10395
rect 1260 10355 1275 10395
rect 1205 10315 1275 10355
rect 1205 10275 1220 10315
rect 1260 10275 1275 10315
rect 1205 10260 1275 10275
rect 1320 12235 1390 12255
rect 1320 12195 1335 12235
rect 1375 12195 1390 12235
rect 1320 12155 1390 12195
rect 1320 12115 1335 12155
rect 1375 12115 1390 12155
rect 1320 12075 1390 12115
rect 1320 12035 1335 12075
rect 1375 12035 1390 12075
rect 1320 11995 1390 12035
rect 1320 11955 1335 11995
rect 1375 11955 1390 11995
rect 1320 11915 1390 11955
rect 1320 11875 1335 11915
rect 1375 11875 1390 11915
rect 1320 11835 1390 11875
rect 1320 11795 1335 11835
rect 1375 11795 1390 11835
rect 1320 11755 1390 11795
rect 1320 11715 1335 11755
rect 1375 11715 1390 11755
rect 1320 11675 1390 11715
rect 1320 11635 1335 11675
rect 1375 11635 1390 11675
rect 1320 11595 1390 11635
rect 1320 11555 1335 11595
rect 1375 11555 1390 11595
rect 1320 11515 1390 11555
rect 1320 11475 1335 11515
rect 1375 11475 1390 11515
rect 1320 11435 1390 11475
rect 1320 11395 1335 11435
rect 1375 11395 1390 11435
rect 1320 11355 1390 11395
rect 1320 11315 1335 11355
rect 1375 11315 1390 11355
rect 1320 11275 1390 11315
rect 1320 11235 1335 11275
rect 1375 11235 1390 11275
rect 1320 11195 1390 11235
rect 1320 11155 1335 11195
rect 1375 11155 1390 11195
rect 1320 11115 1390 11155
rect 1320 11075 1335 11115
rect 1375 11075 1390 11115
rect 1320 11035 1390 11075
rect 1320 10995 1335 11035
rect 1375 10995 1390 11035
rect 1320 10955 1390 10995
rect 1320 10915 1335 10955
rect 1375 10915 1390 10955
rect 1320 10875 1390 10915
rect 1320 10835 1335 10875
rect 1375 10835 1390 10875
rect 1320 10795 1390 10835
rect 1320 10755 1335 10795
rect 1375 10755 1390 10795
rect 1320 10715 1390 10755
rect 1320 10675 1335 10715
rect 1375 10675 1390 10715
rect 1320 10635 1390 10675
rect 1320 10595 1335 10635
rect 1375 10595 1390 10635
rect 1320 10555 1390 10595
rect 1320 10515 1335 10555
rect 1375 10515 1390 10555
rect 1320 10475 1390 10515
rect 1320 10435 1335 10475
rect 1375 10435 1390 10475
rect 1320 10395 1390 10435
rect 1320 10355 1335 10395
rect 1375 10355 1390 10395
rect 1320 10315 1390 10355
rect 1320 10275 1335 10315
rect 1375 10275 1390 10315
rect 1320 10260 1390 10275
rect 1435 12235 1505 12255
rect 1435 12195 1450 12235
rect 1490 12195 1505 12235
rect 1435 12155 1505 12195
rect 1435 12115 1450 12155
rect 1490 12115 1505 12155
rect 1435 12075 1505 12115
rect 1435 12035 1450 12075
rect 1490 12035 1505 12075
rect 1435 11995 1505 12035
rect 1435 11955 1450 11995
rect 1490 11955 1505 11995
rect 1435 11915 1505 11955
rect 1435 11875 1450 11915
rect 1490 11875 1505 11915
rect 1435 11835 1505 11875
rect 1435 11795 1450 11835
rect 1490 11795 1505 11835
rect 1435 11755 1505 11795
rect 1435 11715 1450 11755
rect 1490 11715 1505 11755
rect 1435 11675 1505 11715
rect 1435 11635 1450 11675
rect 1490 11635 1505 11675
rect 1435 11595 1505 11635
rect 1435 11555 1450 11595
rect 1490 11555 1505 11595
rect 1435 11515 1505 11555
rect 1435 11475 1450 11515
rect 1490 11475 1505 11515
rect 1435 11435 1505 11475
rect 1435 11395 1450 11435
rect 1490 11395 1505 11435
rect 1435 11355 1505 11395
rect 1435 11315 1450 11355
rect 1490 11315 1505 11355
rect 1435 11275 1505 11315
rect 1435 11235 1450 11275
rect 1490 11235 1505 11275
rect 1435 11195 1505 11235
rect 1435 11155 1450 11195
rect 1490 11155 1505 11195
rect 1435 11115 1505 11155
rect 1435 11075 1450 11115
rect 1490 11075 1505 11115
rect 1435 11035 1505 11075
rect 1435 10995 1450 11035
rect 1490 10995 1505 11035
rect 1435 10955 1505 10995
rect 1435 10915 1450 10955
rect 1490 10915 1505 10955
rect 1435 10875 1505 10915
rect 1435 10835 1450 10875
rect 1490 10835 1505 10875
rect 1435 10795 1505 10835
rect 1435 10755 1450 10795
rect 1490 10755 1505 10795
rect 1435 10715 1505 10755
rect 1435 10675 1450 10715
rect 1490 10675 1505 10715
rect 1435 10635 1505 10675
rect 1435 10595 1450 10635
rect 1490 10595 1505 10635
rect 1435 10555 1505 10595
rect 1435 10515 1450 10555
rect 1490 10515 1505 10555
rect 1435 10475 1505 10515
rect 1435 10435 1450 10475
rect 1490 10435 1505 10475
rect 1435 10395 1505 10435
rect 1435 10355 1450 10395
rect 1490 10355 1505 10395
rect 1435 10315 1505 10355
rect 1435 10275 1450 10315
rect 1490 10275 1505 10315
rect 1435 10260 1505 10275
rect 1550 12235 1620 12255
rect 1550 12195 1565 12235
rect 1605 12195 1620 12235
rect 1550 12155 1620 12195
rect 1550 12115 1565 12155
rect 1605 12115 1620 12155
rect 1550 12075 1620 12115
rect 1550 12035 1565 12075
rect 1605 12035 1620 12075
rect 1550 11995 1620 12035
rect 1550 11955 1565 11995
rect 1605 11955 1620 11995
rect 1550 11915 1620 11955
rect 1550 11875 1565 11915
rect 1605 11875 1620 11915
rect 1550 11835 1620 11875
rect 1550 11795 1565 11835
rect 1605 11795 1620 11835
rect 1550 11755 1620 11795
rect 1550 11715 1565 11755
rect 1605 11715 1620 11755
rect 1550 11675 1620 11715
rect 1550 11635 1565 11675
rect 1605 11635 1620 11675
rect 1550 11595 1620 11635
rect 1550 11555 1565 11595
rect 1605 11555 1620 11595
rect 1550 11515 1620 11555
rect 1550 11475 1565 11515
rect 1605 11475 1620 11515
rect 1550 11435 1620 11475
rect 1550 11395 1565 11435
rect 1605 11395 1620 11435
rect 1550 11355 1620 11395
rect 1550 11315 1565 11355
rect 1605 11315 1620 11355
rect 1550 11275 1620 11315
rect 1550 11235 1565 11275
rect 1605 11235 1620 11275
rect 1550 11195 1620 11235
rect 1550 11155 1565 11195
rect 1605 11155 1620 11195
rect 1550 11115 1620 11155
rect 1550 11075 1565 11115
rect 1605 11075 1620 11115
rect 1550 11035 1620 11075
rect 1550 10995 1565 11035
rect 1605 10995 1620 11035
rect 1550 10955 1620 10995
rect 1550 10915 1565 10955
rect 1605 10915 1620 10955
rect 1550 10875 1620 10915
rect 1550 10835 1565 10875
rect 1605 10835 1620 10875
rect 1550 10795 1620 10835
rect 1550 10755 1565 10795
rect 1605 10755 1620 10795
rect 1550 10715 1620 10755
rect 1550 10675 1565 10715
rect 1605 10675 1620 10715
rect 1550 10635 1620 10675
rect 1550 10595 1565 10635
rect 1605 10595 1620 10635
rect 1550 10555 1620 10595
rect 1550 10515 1565 10555
rect 1605 10515 1620 10555
rect 1550 10475 1620 10515
rect 1550 10435 1565 10475
rect 1605 10435 1620 10475
rect 1550 10395 1620 10435
rect 1550 10355 1565 10395
rect 1605 10355 1620 10395
rect 1550 10315 1620 10355
rect 1550 10275 1565 10315
rect 1605 10275 1620 10315
rect 1550 10260 1620 10275
rect 1665 12235 1735 12255
rect 1665 12195 1680 12235
rect 1720 12195 1735 12235
rect 1665 12155 1735 12195
rect 1665 12115 1680 12155
rect 1720 12115 1735 12155
rect 1665 12075 1735 12115
rect 1665 12035 1680 12075
rect 1720 12035 1735 12075
rect 1665 11995 1735 12035
rect 1665 11955 1680 11995
rect 1720 11955 1735 11995
rect 1665 11915 1735 11955
rect 1665 11875 1680 11915
rect 1720 11875 1735 11915
rect 1665 11835 1735 11875
rect 1665 11795 1680 11835
rect 1720 11795 1735 11835
rect 1665 11755 1735 11795
rect 1665 11715 1680 11755
rect 1720 11715 1735 11755
rect 1665 11675 1735 11715
rect 1665 11635 1680 11675
rect 1720 11635 1735 11675
rect 1665 11595 1735 11635
rect 1665 11555 1680 11595
rect 1720 11555 1735 11595
rect 1665 11515 1735 11555
rect 1665 11475 1680 11515
rect 1720 11475 1735 11515
rect 1665 11435 1735 11475
rect 1665 11395 1680 11435
rect 1720 11395 1735 11435
rect 1665 11355 1735 11395
rect 1665 11315 1680 11355
rect 1720 11315 1735 11355
rect 1665 11275 1735 11315
rect 1665 11235 1680 11275
rect 1720 11235 1735 11275
rect 1665 11195 1735 11235
rect 1665 11155 1680 11195
rect 1720 11155 1735 11195
rect 1665 11115 1735 11155
rect 1665 11075 1680 11115
rect 1720 11075 1735 11115
rect 1665 11035 1735 11075
rect 1665 10995 1680 11035
rect 1720 10995 1735 11035
rect 1665 10955 1735 10995
rect 1665 10915 1680 10955
rect 1720 10915 1735 10955
rect 1665 10875 1735 10915
rect 1665 10835 1680 10875
rect 1720 10835 1735 10875
rect 1665 10795 1735 10835
rect 1665 10755 1680 10795
rect 1720 10755 1735 10795
rect 1665 10715 1735 10755
rect 1665 10675 1680 10715
rect 1720 10675 1735 10715
rect 1665 10635 1735 10675
rect 1665 10595 1680 10635
rect 1720 10595 1735 10635
rect 1665 10555 1735 10595
rect 1665 10515 1680 10555
rect 1720 10515 1735 10555
rect 1665 10475 1735 10515
rect 1665 10435 1680 10475
rect 1720 10435 1735 10475
rect 1665 10395 1735 10435
rect 1665 10355 1680 10395
rect 1720 10355 1735 10395
rect 1665 10315 1735 10355
rect 1665 10275 1680 10315
rect 1720 10275 1735 10315
rect 1665 10260 1735 10275
rect 1780 12235 1850 12255
rect 1780 12195 1795 12235
rect 1835 12195 1850 12235
rect 1780 12155 1850 12195
rect 1780 12115 1795 12155
rect 1835 12115 1850 12155
rect 1780 12075 1850 12115
rect 1780 12035 1795 12075
rect 1835 12035 1850 12075
rect 1780 11995 1850 12035
rect 1780 11955 1795 11995
rect 1835 11955 1850 11995
rect 1780 11915 1850 11955
rect 1780 11875 1795 11915
rect 1835 11875 1850 11915
rect 1780 11835 1850 11875
rect 1780 11795 1795 11835
rect 1835 11795 1850 11835
rect 1780 11755 1850 11795
rect 1780 11715 1795 11755
rect 1835 11715 1850 11755
rect 1780 11675 1850 11715
rect 1780 11635 1795 11675
rect 1835 11635 1850 11675
rect 1780 11595 1850 11635
rect 1780 11555 1795 11595
rect 1835 11555 1850 11595
rect 1780 11515 1850 11555
rect 1780 11475 1795 11515
rect 1835 11475 1850 11515
rect 1780 11435 1850 11475
rect 1780 11395 1795 11435
rect 1835 11395 1850 11435
rect 1780 11355 1850 11395
rect 1780 11315 1795 11355
rect 1835 11315 1850 11355
rect 1780 11275 1850 11315
rect 1780 11235 1795 11275
rect 1835 11235 1850 11275
rect 1780 11195 1850 11235
rect 1780 11155 1795 11195
rect 1835 11155 1850 11195
rect 1780 11115 1850 11155
rect 1780 11075 1795 11115
rect 1835 11075 1850 11115
rect 1780 11035 1850 11075
rect 1780 10995 1795 11035
rect 1835 10995 1850 11035
rect 1780 10955 1850 10995
rect 1780 10915 1795 10955
rect 1835 10915 1850 10955
rect 1780 10875 1850 10915
rect 1780 10835 1795 10875
rect 1835 10835 1850 10875
rect 1780 10795 1850 10835
rect 1780 10755 1795 10795
rect 1835 10755 1850 10795
rect 1780 10715 1850 10755
rect 1780 10675 1795 10715
rect 1835 10675 1850 10715
rect 1780 10635 1850 10675
rect 1780 10595 1795 10635
rect 1835 10595 1850 10635
rect 1780 10555 1850 10595
rect 1780 10515 1795 10555
rect 1835 10515 1850 10555
rect 1780 10475 1850 10515
rect 1780 10435 1795 10475
rect 1835 10435 1850 10475
rect 1780 10395 1850 10435
rect 1780 10355 1795 10395
rect 1835 10355 1850 10395
rect 1780 10315 1850 10355
rect 1780 10275 1795 10315
rect 1835 10275 1850 10315
rect 1780 10260 1850 10275
rect 1895 12235 1965 12255
rect 1895 12195 1910 12235
rect 1950 12195 1965 12235
rect 1895 12155 1965 12195
rect 1895 12115 1910 12155
rect 1950 12115 1965 12155
rect 1895 12075 1965 12115
rect 1895 12035 1910 12075
rect 1950 12035 1965 12075
rect 1895 11995 1965 12035
rect 1895 11955 1910 11995
rect 1950 11955 1965 11995
rect 1895 11915 1965 11955
rect 1895 11875 1910 11915
rect 1950 11875 1965 11915
rect 1895 11835 1965 11875
rect 1895 11795 1910 11835
rect 1950 11795 1965 11835
rect 1895 11755 1965 11795
rect 1895 11715 1910 11755
rect 1950 11715 1965 11755
rect 1895 11675 1965 11715
rect 1895 11635 1910 11675
rect 1950 11635 1965 11675
rect 1895 11595 1965 11635
rect 1895 11555 1910 11595
rect 1950 11555 1965 11595
rect 1895 11515 1965 11555
rect 1895 11475 1910 11515
rect 1950 11475 1965 11515
rect 1895 11435 1965 11475
rect 1895 11395 1910 11435
rect 1950 11395 1965 11435
rect 1895 11355 1965 11395
rect 1895 11315 1910 11355
rect 1950 11315 1965 11355
rect 1895 11275 1965 11315
rect 1895 11235 1910 11275
rect 1950 11235 1965 11275
rect 1895 11195 1965 11235
rect 1895 11155 1910 11195
rect 1950 11155 1965 11195
rect 1895 11115 1965 11155
rect 1895 11075 1910 11115
rect 1950 11075 1965 11115
rect 1895 11035 1965 11075
rect 1895 10995 1910 11035
rect 1950 10995 1965 11035
rect 1895 10955 1965 10995
rect 1895 10915 1910 10955
rect 1950 10915 1965 10955
rect 1895 10875 1965 10915
rect 1895 10835 1910 10875
rect 1950 10835 1965 10875
rect 1895 10795 1965 10835
rect 1895 10755 1910 10795
rect 1950 10755 1965 10795
rect 1895 10715 1965 10755
rect 1895 10675 1910 10715
rect 1950 10675 1965 10715
rect 1895 10635 1965 10675
rect 1895 10595 1910 10635
rect 1950 10595 1965 10635
rect 1895 10555 1965 10595
rect 1895 10515 1910 10555
rect 1950 10515 1965 10555
rect 1895 10475 1965 10515
rect 1895 10435 1910 10475
rect 1950 10435 1965 10475
rect 1895 10395 1965 10435
rect 1895 10355 1910 10395
rect 1950 10355 1965 10395
rect 1895 10315 1965 10355
rect 1895 10275 1910 10315
rect 1950 10275 1965 10315
rect 1895 10260 1965 10275
rect 2010 12235 2080 12255
rect 2010 12195 2025 12235
rect 2065 12195 2080 12235
rect 2010 12155 2080 12195
rect 2010 12115 2025 12155
rect 2065 12115 2080 12155
rect 2010 12075 2080 12115
rect 2010 12035 2025 12075
rect 2065 12035 2080 12075
rect 2010 11995 2080 12035
rect 2010 11955 2025 11995
rect 2065 11955 2080 11995
rect 2010 11915 2080 11955
rect 2010 11875 2025 11915
rect 2065 11875 2080 11915
rect 2010 11835 2080 11875
rect 2010 11795 2025 11835
rect 2065 11795 2080 11835
rect 2010 11755 2080 11795
rect 2010 11715 2025 11755
rect 2065 11715 2080 11755
rect 2010 11675 2080 11715
rect 2010 11635 2025 11675
rect 2065 11635 2080 11675
rect 2010 11595 2080 11635
rect 2010 11555 2025 11595
rect 2065 11555 2080 11595
rect 2010 11515 2080 11555
rect 2010 11475 2025 11515
rect 2065 11475 2080 11515
rect 2010 11435 2080 11475
rect 2010 11395 2025 11435
rect 2065 11395 2080 11435
rect 2010 11355 2080 11395
rect 2010 11315 2025 11355
rect 2065 11315 2080 11355
rect 2010 11275 2080 11315
rect 2010 11235 2025 11275
rect 2065 11235 2080 11275
rect 2010 11195 2080 11235
rect 2010 11155 2025 11195
rect 2065 11155 2080 11195
rect 2010 11115 2080 11155
rect 2010 11075 2025 11115
rect 2065 11075 2080 11115
rect 2010 11035 2080 11075
rect 2010 10995 2025 11035
rect 2065 10995 2080 11035
rect 2010 10955 2080 10995
rect 2010 10915 2025 10955
rect 2065 10915 2080 10955
rect 2010 10875 2080 10915
rect 2010 10835 2025 10875
rect 2065 10835 2080 10875
rect 2010 10795 2080 10835
rect 2010 10755 2025 10795
rect 2065 10755 2080 10795
rect 2010 10715 2080 10755
rect 2010 10675 2025 10715
rect 2065 10675 2080 10715
rect 2010 10635 2080 10675
rect 2010 10595 2025 10635
rect 2065 10595 2080 10635
rect 2010 10555 2080 10595
rect 2010 10515 2025 10555
rect 2065 10515 2080 10555
rect 2010 10475 2080 10515
rect 2010 10435 2025 10475
rect 2065 10435 2080 10475
rect 2010 10395 2080 10435
rect 2010 10355 2025 10395
rect 2065 10355 2080 10395
rect 2010 10315 2080 10355
rect 2010 10275 2025 10315
rect 2065 10275 2080 10315
rect 2010 10260 2080 10275
rect 2125 12235 2195 12255
rect 2125 12195 2140 12235
rect 2180 12195 2195 12235
rect 2125 12155 2195 12195
rect 2125 12115 2140 12155
rect 2180 12115 2195 12155
rect 2125 12075 2195 12115
rect 2125 12035 2140 12075
rect 2180 12035 2195 12075
rect 2125 11995 2195 12035
rect 2125 11955 2140 11995
rect 2180 11955 2195 11995
rect 2125 11915 2195 11955
rect 2125 11875 2140 11915
rect 2180 11875 2195 11915
rect 2125 11835 2195 11875
rect 2125 11795 2140 11835
rect 2180 11795 2195 11835
rect 2125 11755 2195 11795
rect 2125 11715 2140 11755
rect 2180 11715 2195 11755
rect 2125 11675 2195 11715
rect 2125 11635 2140 11675
rect 2180 11635 2195 11675
rect 2125 11595 2195 11635
rect 2125 11555 2140 11595
rect 2180 11555 2195 11595
rect 2125 11515 2195 11555
rect 2125 11475 2140 11515
rect 2180 11475 2195 11515
rect 2125 11435 2195 11475
rect 2125 11395 2140 11435
rect 2180 11395 2195 11435
rect 2125 11355 2195 11395
rect 2125 11315 2140 11355
rect 2180 11315 2195 11355
rect 2125 11275 2195 11315
rect 2125 11235 2140 11275
rect 2180 11235 2195 11275
rect 2125 11195 2195 11235
rect 2125 11155 2140 11195
rect 2180 11155 2195 11195
rect 2125 11115 2195 11155
rect 2125 11075 2140 11115
rect 2180 11075 2195 11115
rect 2125 11035 2195 11075
rect 2125 10995 2140 11035
rect 2180 10995 2195 11035
rect 2125 10955 2195 10995
rect 2125 10915 2140 10955
rect 2180 10915 2195 10955
rect 2125 10875 2195 10915
rect 2125 10835 2140 10875
rect 2180 10835 2195 10875
rect 2125 10795 2195 10835
rect 2125 10755 2140 10795
rect 2180 10755 2195 10795
rect 2125 10715 2195 10755
rect 2125 10675 2140 10715
rect 2180 10675 2195 10715
rect 2125 10635 2195 10675
rect 2125 10595 2140 10635
rect 2180 10595 2195 10635
rect 2125 10555 2195 10595
rect 2125 10515 2140 10555
rect 2180 10515 2195 10555
rect 2125 10475 2195 10515
rect 2125 10435 2140 10475
rect 2180 10435 2195 10475
rect 2125 10395 2195 10435
rect 2125 10355 2140 10395
rect 2180 10355 2195 10395
rect 2125 10315 2195 10355
rect 2125 10275 2140 10315
rect 2180 10275 2195 10315
rect 2125 10260 2195 10275
rect 2240 12235 2310 12255
rect 2240 12195 2255 12235
rect 2295 12195 2310 12235
rect 2240 12155 2310 12195
rect 2240 12115 2255 12155
rect 2295 12115 2310 12155
rect 2240 12075 2310 12115
rect 2240 12035 2255 12075
rect 2295 12035 2310 12075
rect 2240 11995 2310 12035
rect 2240 11955 2255 11995
rect 2295 11955 2310 11995
rect 2240 11915 2310 11955
rect 2240 11875 2255 11915
rect 2295 11875 2310 11915
rect 2240 11835 2310 11875
rect 2240 11795 2255 11835
rect 2295 11795 2310 11835
rect 2240 11755 2310 11795
rect 2240 11715 2255 11755
rect 2295 11715 2310 11755
rect 2240 11675 2310 11715
rect 2240 11635 2255 11675
rect 2295 11635 2310 11675
rect 2240 11595 2310 11635
rect 2240 11555 2255 11595
rect 2295 11555 2310 11595
rect 2240 11515 2310 11555
rect 2240 11475 2255 11515
rect 2295 11475 2310 11515
rect 2240 11435 2310 11475
rect 2240 11395 2255 11435
rect 2295 11395 2310 11435
rect 2240 11355 2310 11395
rect 2240 11315 2255 11355
rect 2295 11315 2310 11355
rect 2240 11275 2310 11315
rect 2240 11235 2255 11275
rect 2295 11235 2310 11275
rect 2240 11195 2310 11235
rect 2240 11155 2255 11195
rect 2295 11155 2310 11195
rect 2240 11115 2310 11155
rect 2240 11075 2255 11115
rect 2295 11075 2310 11115
rect 2240 11035 2310 11075
rect 2240 10995 2255 11035
rect 2295 10995 2310 11035
rect 2240 10955 2310 10995
rect 2240 10915 2255 10955
rect 2295 10915 2310 10955
rect 2240 10875 2310 10915
rect 2240 10835 2255 10875
rect 2295 10835 2310 10875
rect 2240 10795 2310 10835
rect 2240 10755 2255 10795
rect 2295 10755 2310 10795
rect 2240 10715 2310 10755
rect 2240 10675 2255 10715
rect 2295 10675 2310 10715
rect 2240 10635 2310 10675
rect 2240 10595 2255 10635
rect 2295 10595 2310 10635
rect 2240 10555 2310 10595
rect 2240 10515 2255 10555
rect 2295 10515 2310 10555
rect 2240 10475 2310 10515
rect 2240 10435 2255 10475
rect 2295 10435 2310 10475
rect 2240 10395 2310 10435
rect 2240 10355 2255 10395
rect 2295 10355 2310 10395
rect 2240 10315 2310 10355
rect 2240 10275 2255 10315
rect 2295 10275 2310 10315
rect 2240 10260 2310 10275
rect 2355 12235 2425 12255
rect 2355 12195 2370 12235
rect 2410 12195 2425 12235
rect 2355 12155 2425 12195
rect 2355 12115 2370 12155
rect 2410 12115 2425 12155
rect 2355 12075 2425 12115
rect 2355 12035 2370 12075
rect 2410 12035 2425 12075
rect 2355 11995 2425 12035
rect 2355 11955 2370 11995
rect 2410 11955 2425 11995
rect 2355 11915 2425 11955
rect 2355 11875 2370 11915
rect 2410 11875 2425 11915
rect 2355 11835 2425 11875
rect 2355 11795 2370 11835
rect 2410 11795 2425 11835
rect 2355 11755 2425 11795
rect 2355 11715 2370 11755
rect 2410 11715 2425 11755
rect 2355 11675 2425 11715
rect 2355 11635 2370 11675
rect 2410 11635 2425 11675
rect 2355 11595 2425 11635
rect 2355 11555 2370 11595
rect 2410 11555 2425 11595
rect 2355 11515 2425 11555
rect 2355 11475 2370 11515
rect 2410 11475 2425 11515
rect 2355 11435 2425 11475
rect 2355 11395 2370 11435
rect 2410 11395 2425 11435
rect 2355 11355 2425 11395
rect 2355 11315 2370 11355
rect 2410 11315 2425 11355
rect 2355 11275 2425 11315
rect 2355 11235 2370 11275
rect 2410 11235 2425 11275
rect 2355 11195 2425 11235
rect 2355 11155 2370 11195
rect 2410 11155 2425 11195
rect 2355 11115 2425 11155
rect 2355 11075 2370 11115
rect 2410 11075 2425 11115
rect 2355 11035 2425 11075
rect 2355 10995 2370 11035
rect 2410 10995 2425 11035
rect 2355 10955 2425 10995
rect 2355 10915 2370 10955
rect 2410 10915 2425 10955
rect 2355 10875 2425 10915
rect 2355 10835 2370 10875
rect 2410 10835 2425 10875
rect 2355 10795 2425 10835
rect 2355 10755 2370 10795
rect 2410 10755 2425 10795
rect 2355 10715 2425 10755
rect 2355 10675 2370 10715
rect 2410 10675 2425 10715
rect 2355 10635 2425 10675
rect 2355 10595 2370 10635
rect 2410 10595 2425 10635
rect 2355 10555 2425 10595
rect 2355 10515 2370 10555
rect 2410 10515 2425 10555
rect 2355 10475 2425 10515
rect 2355 10435 2370 10475
rect 2410 10435 2425 10475
rect 2355 10395 2425 10435
rect 2355 10355 2370 10395
rect 2410 10355 2425 10395
rect 2355 10315 2425 10355
rect 2355 10275 2370 10315
rect 2410 10275 2425 10315
rect 2355 10260 2425 10275
rect 2470 12235 2540 12255
rect 2470 12195 2485 12235
rect 2525 12195 2540 12235
rect 2470 12155 2540 12195
rect 2470 12115 2485 12155
rect 2525 12115 2540 12155
rect 2470 12075 2540 12115
rect 2470 12035 2485 12075
rect 2525 12035 2540 12075
rect 2470 11995 2540 12035
rect 2470 11955 2485 11995
rect 2525 11955 2540 11995
rect 2470 11915 2540 11955
rect 2470 11875 2485 11915
rect 2525 11875 2540 11915
rect 2470 11835 2540 11875
rect 2470 11795 2485 11835
rect 2525 11795 2540 11835
rect 2470 11755 2540 11795
rect 2470 11715 2485 11755
rect 2525 11715 2540 11755
rect 2470 11675 2540 11715
rect 2470 11635 2485 11675
rect 2525 11635 2540 11675
rect 2470 11595 2540 11635
rect 2470 11555 2485 11595
rect 2525 11555 2540 11595
rect 2470 11515 2540 11555
rect 2470 11475 2485 11515
rect 2525 11475 2540 11515
rect 2470 11435 2540 11475
rect 2470 11395 2485 11435
rect 2525 11395 2540 11435
rect 2470 11355 2540 11395
rect 2470 11315 2485 11355
rect 2525 11315 2540 11355
rect 2470 11275 2540 11315
rect 2470 11235 2485 11275
rect 2525 11235 2540 11275
rect 2470 11195 2540 11235
rect 2470 11155 2485 11195
rect 2525 11155 2540 11195
rect 2470 11115 2540 11155
rect 2470 11075 2485 11115
rect 2525 11075 2540 11115
rect 2470 11035 2540 11075
rect 2470 10995 2485 11035
rect 2525 10995 2540 11035
rect 2470 10955 2540 10995
rect 2470 10915 2485 10955
rect 2525 10915 2540 10955
rect 2470 10875 2540 10915
rect 2470 10835 2485 10875
rect 2525 10835 2540 10875
rect 2470 10795 2540 10835
rect 2470 10755 2485 10795
rect 2525 10755 2540 10795
rect 2470 10715 2540 10755
rect 2470 10675 2485 10715
rect 2525 10675 2540 10715
rect 2470 10635 2540 10675
rect 2470 10595 2485 10635
rect 2525 10595 2540 10635
rect 2470 10555 2540 10595
rect 2470 10515 2485 10555
rect 2525 10515 2540 10555
rect 2470 10475 2540 10515
rect 2470 10435 2485 10475
rect 2525 10435 2540 10475
rect 2470 10395 2540 10435
rect 2470 10355 2485 10395
rect 2525 10355 2540 10395
rect 2470 10315 2540 10355
rect 2470 10275 2485 10315
rect 2525 10275 2540 10315
rect 2470 10260 2540 10275
rect 2670 12155 2740 12270
rect 2670 12115 2685 12155
rect 2725 12115 2740 12155
rect 2670 11995 2740 12115
rect 2670 11955 2685 11995
rect 2725 11955 2740 11995
rect 2670 11835 2740 11955
rect 2670 11795 2685 11835
rect 2725 11795 2740 11835
rect 2670 11675 2740 11795
rect 2670 11635 2685 11675
rect 2725 11635 2740 11675
rect 2670 11515 2740 11635
rect 2670 11475 2685 11515
rect 2725 11475 2740 11515
rect 2670 11355 2740 11475
rect 2670 11315 2685 11355
rect 2725 11315 2740 11355
rect 2670 11195 2740 11315
rect 2670 11155 2685 11195
rect 2725 11155 2740 11195
rect 2670 10955 2740 11155
rect 2670 10915 2685 10955
rect 2725 10915 2740 10955
rect 2670 10795 2740 10915
rect 2670 10755 2685 10795
rect 2725 10755 2740 10795
rect 2670 10635 2740 10755
rect 2670 10595 2685 10635
rect 2725 10595 2740 10635
rect 2670 10475 2740 10595
rect 2670 10435 2685 10475
rect 2725 10435 2740 10475
rect 2670 10315 2740 10435
rect 2670 10275 2685 10315
rect 2725 10275 2740 10315
rect 2670 10245 2740 10275
rect -405 10030 865 10045
rect -405 9990 -390 10030
rect -350 9990 -230 10030
rect -190 9990 -70 10030
rect -30 9990 90 10030
rect 130 9990 250 10030
rect 290 9990 410 10030
rect 450 9990 570 10030
rect 610 9990 730 10030
rect 770 9990 865 10030
rect -405 9975 865 9990
rect 1025 10025 1110 10040
rect 1025 9975 1040 10025
rect 1095 9975 1110 10025
rect 1275 10030 2545 10045
rect 1275 9990 1290 10030
rect 1330 9990 1450 10030
rect 1490 9990 1610 10030
rect 1650 9990 1770 10030
rect 1810 9990 1930 10030
rect 1970 9990 2090 10030
rect 2130 9990 2250 10030
rect 2290 9990 2410 10030
rect 2450 9990 2545 10030
rect 1275 9975 2545 9990
rect 1025 9960 1110 9975
<< viali >>
rect -390 12435 -350 12475
rect -230 12435 -190 12475
rect -70 12435 -30 12475
rect 90 12435 130 12475
rect 250 12435 290 12475
rect 410 12435 450 12475
rect 570 12435 610 12475
rect 730 12435 770 12475
rect 1290 12435 1330 12475
rect 1450 12435 1490 12475
rect 1610 12435 1650 12475
rect 1770 12435 1810 12475
rect 1930 12435 1970 12475
rect 2090 12435 2130 12475
rect 2250 12435 2290 12475
rect 2410 12435 2450 12475
rect -590 12195 -550 12235
rect -590 12035 -550 12075
rect -590 11875 -550 11915
rect -590 11715 -550 11755
rect -590 11555 -550 11595
rect -590 11395 -550 11435
rect -590 11235 -550 11275
rect -590 11075 -550 11115
rect -590 10915 -550 10955
rect -590 10755 -550 10795
rect -590 10595 -550 10635
rect -590 10435 -550 10475
rect -590 10275 -550 10315
rect -390 12195 -350 12235
rect -390 12115 -350 12155
rect -390 12035 -350 12075
rect -390 11955 -350 11995
rect -390 11875 -350 11915
rect -390 11795 -350 11835
rect -390 11715 -350 11755
rect -390 11635 -350 11675
rect -390 11555 -350 11595
rect -390 11475 -350 11515
rect -390 11395 -350 11435
rect -390 11315 -350 11355
rect -390 11235 -350 11275
rect -390 11155 -350 11195
rect -390 11075 -350 11115
rect -390 10995 -350 11035
rect -390 10915 -350 10955
rect -390 10835 -350 10875
rect -390 10755 -350 10795
rect -390 10675 -350 10715
rect -390 10595 -350 10635
rect -390 10515 -350 10555
rect -390 10435 -350 10475
rect -390 10355 -350 10395
rect -390 10275 -350 10315
rect -275 12195 -235 12235
rect -275 12115 -235 12155
rect -275 12035 -235 12075
rect -275 11955 -235 11995
rect -275 11875 -235 11915
rect -275 11795 -235 11835
rect -275 11715 -235 11755
rect -275 11635 -235 11675
rect -275 11555 -235 11595
rect -275 11475 -235 11515
rect -275 11395 -235 11435
rect -275 11315 -235 11355
rect -275 11235 -235 11275
rect -275 11155 -235 11195
rect -275 11075 -235 11115
rect -275 10995 -235 11035
rect -275 10915 -235 10955
rect -275 10835 -235 10875
rect -275 10755 -235 10795
rect -275 10675 -235 10715
rect -275 10595 -235 10635
rect -275 10515 -235 10555
rect -275 10435 -235 10475
rect -275 10355 -235 10395
rect -275 10275 -235 10315
rect -160 12195 -120 12235
rect -160 12115 -120 12155
rect -160 12035 -120 12075
rect -160 11955 -120 11995
rect -160 11875 -120 11915
rect -160 11795 -120 11835
rect -160 11715 -120 11755
rect -160 11635 -120 11675
rect -160 11555 -120 11595
rect -160 11475 -120 11515
rect -160 11395 -120 11435
rect -160 11315 -120 11355
rect -160 11235 -120 11275
rect -160 11155 -120 11195
rect -160 11075 -120 11115
rect -160 10995 -120 11035
rect -160 10915 -120 10955
rect -160 10835 -120 10875
rect -160 10755 -120 10795
rect -160 10675 -120 10715
rect -160 10595 -120 10635
rect -160 10515 -120 10555
rect -160 10435 -120 10475
rect -160 10355 -120 10395
rect -160 10275 -120 10315
rect -45 12195 -5 12235
rect -45 12115 -5 12155
rect -45 12035 -5 12075
rect -45 11955 -5 11995
rect -45 11875 -5 11915
rect -45 11795 -5 11835
rect -45 11715 -5 11755
rect -45 11635 -5 11675
rect -45 11555 -5 11595
rect -45 11475 -5 11515
rect -45 11395 -5 11435
rect -45 11315 -5 11355
rect -45 11235 -5 11275
rect -45 11155 -5 11195
rect -45 11075 -5 11115
rect -45 10995 -5 11035
rect -45 10915 -5 10955
rect -45 10835 -5 10875
rect -45 10755 -5 10795
rect -45 10675 -5 10715
rect -45 10595 -5 10635
rect -45 10515 -5 10555
rect -45 10435 -5 10475
rect -45 10355 -5 10395
rect -45 10275 -5 10315
rect 70 12195 110 12235
rect 70 12115 110 12155
rect 70 12035 110 12075
rect 70 11955 110 11995
rect 70 11875 110 11915
rect 70 11795 110 11835
rect 70 11715 110 11755
rect 70 11635 110 11675
rect 70 11555 110 11595
rect 70 11475 110 11515
rect 70 11395 110 11435
rect 70 11315 110 11355
rect 70 11235 110 11275
rect 70 11155 110 11195
rect 70 11075 110 11115
rect 70 10995 110 11035
rect 70 10915 110 10955
rect 70 10835 110 10875
rect 70 10755 110 10795
rect 70 10675 110 10715
rect 70 10595 110 10635
rect 70 10515 110 10555
rect 70 10435 110 10475
rect 70 10355 110 10395
rect 70 10275 110 10315
rect 185 12195 225 12235
rect 185 12115 225 12155
rect 185 12035 225 12075
rect 185 11955 225 11995
rect 185 11875 225 11915
rect 185 11795 225 11835
rect 185 11715 225 11755
rect 185 11635 225 11675
rect 185 11555 225 11595
rect 185 11475 225 11515
rect 185 11395 225 11435
rect 185 11315 225 11355
rect 185 11235 225 11275
rect 185 11155 225 11195
rect 185 11075 225 11115
rect 185 10995 225 11035
rect 185 10915 225 10955
rect 185 10835 225 10875
rect 185 10755 225 10795
rect 185 10675 225 10715
rect 185 10595 225 10635
rect 185 10515 225 10555
rect 185 10435 225 10475
rect 185 10355 225 10395
rect 185 10275 225 10315
rect 300 12195 340 12235
rect 300 12115 340 12155
rect 300 12035 340 12075
rect 300 11955 340 11995
rect 300 11875 340 11915
rect 300 11795 340 11835
rect 300 11715 340 11755
rect 300 11635 340 11675
rect 300 11555 340 11595
rect 300 11475 340 11515
rect 300 11395 340 11435
rect 300 11315 340 11355
rect 300 11235 340 11275
rect 300 11155 340 11195
rect 300 11075 340 11115
rect 300 10995 340 11035
rect 300 10915 340 10955
rect 300 10835 340 10875
rect 300 10755 340 10795
rect 300 10675 340 10715
rect 300 10595 340 10635
rect 300 10515 340 10555
rect 300 10435 340 10475
rect 300 10355 340 10395
rect 300 10275 340 10315
rect 415 12195 455 12235
rect 415 12115 455 12155
rect 415 12035 455 12075
rect 415 11955 455 11995
rect 415 11875 455 11915
rect 415 11795 455 11835
rect 415 11715 455 11755
rect 415 11635 455 11675
rect 415 11555 455 11595
rect 415 11475 455 11515
rect 415 11395 455 11435
rect 415 11315 455 11355
rect 415 11235 455 11275
rect 415 11155 455 11195
rect 415 11075 455 11115
rect 415 10995 455 11035
rect 415 10915 455 10955
rect 415 10835 455 10875
rect 415 10755 455 10795
rect 415 10675 455 10715
rect 415 10595 455 10635
rect 415 10515 455 10555
rect 415 10435 455 10475
rect 415 10355 455 10395
rect 415 10275 455 10315
rect 530 12195 570 12235
rect 530 12115 570 12155
rect 530 12035 570 12075
rect 530 11955 570 11995
rect 530 11875 570 11915
rect 530 11795 570 11835
rect 530 11715 570 11755
rect 530 11635 570 11675
rect 530 11555 570 11595
rect 530 11475 570 11515
rect 530 11395 570 11435
rect 530 11315 570 11355
rect 530 11235 570 11275
rect 530 11155 570 11195
rect 530 11075 570 11115
rect 530 10995 570 11035
rect 530 10915 570 10955
rect 530 10835 570 10875
rect 530 10755 570 10795
rect 530 10675 570 10715
rect 530 10595 570 10635
rect 530 10515 570 10555
rect 530 10435 570 10475
rect 530 10355 570 10395
rect 530 10275 570 10315
rect 645 12195 685 12235
rect 645 12115 685 12155
rect 645 12035 685 12075
rect 645 11955 685 11995
rect 645 11875 685 11915
rect 645 11795 685 11835
rect 645 11715 685 11755
rect 645 11635 685 11675
rect 645 11555 685 11595
rect 645 11475 685 11515
rect 645 11395 685 11435
rect 645 11315 685 11355
rect 645 11235 685 11275
rect 645 11155 685 11195
rect 645 11075 685 11115
rect 645 10995 685 11035
rect 645 10915 685 10955
rect 645 10835 685 10875
rect 645 10755 685 10795
rect 645 10675 685 10715
rect 645 10595 685 10635
rect 645 10515 685 10555
rect 645 10435 685 10475
rect 645 10355 685 10395
rect 645 10275 685 10315
rect 760 12195 800 12235
rect 760 12115 800 12155
rect 760 12035 800 12075
rect 760 11955 800 11995
rect 760 11875 800 11915
rect 760 11795 800 11835
rect 760 11715 800 11755
rect 760 11635 800 11675
rect 760 11555 800 11595
rect 760 11475 800 11515
rect 760 11395 800 11435
rect 760 11315 800 11355
rect 760 11235 800 11275
rect 760 11155 800 11195
rect 760 11075 800 11115
rect 760 10995 800 11035
rect 760 10915 800 10955
rect 760 10835 800 10875
rect 760 10755 800 10795
rect 760 10675 800 10715
rect 760 10595 800 10635
rect 760 10515 800 10555
rect 760 10435 800 10475
rect 760 10355 800 10395
rect 760 10275 800 10315
rect 875 12195 915 12235
rect 875 12115 915 12155
rect 875 12035 915 12075
rect 875 11955 915 11995
rect 875 11875 915 11915
rect 875 11795 915 11835
rect 875 11715 915 11755
rect 875 11635 915 11675
rect 875 11555 915 11595
rect 875 11475 915 11515
rect 875 11395 915 11435
rect 875 11315 915 11355
rect 875 11235 915 11275
rect 875 11155 915 11195
rect 875 11075 915 11115
rect 875 10995 915 11035
rect 875 10915 915 10955
rect 875 10835 915 10875
rect 875 10755 915 10795
rect 875 10675 915 10715
rect 875 10595 915 10635
rect 875 10515 915 10555
rect 875 10435 915 10475
rect 875 10355 915 10395
rect 875 10275 915 10315
rect 990 12195 1030 12235
rect 990 12115 1030 12155
rect 990 12035 1030 12075
rect 990 11955 1030 11995
rect 990 11875 1030 11915
rect 990 11795 1030 11835
rect 990 11715 1030 11755
rect 990 11635 1030 11675
rect 990 11555 1030 11595
rect 990 11475 1030 11515
rect 990 11395 1030 11435
rect 990 11315 1030 11355
rect 990 11235 1030 11275
rect 990 11155 1030 11195
rect 990 11075 1030 11115
rect 990 10995 1030 11035
rect 990 10915 1030 10955
rect 990 10835 1030 10875
rect 990 10755 1030 10795
rect 990 10675 1030 10715
rect 990 10595 1030 10635
rect 990 10515 1030 10555
rect 990 10435 1030 10475
rect 990 10355 1030 10395
rect 990 10275 1030 10315
rect 1105 12195 1145 12235
rect 1105 12115 1145 12155
rect 1105 12035 1145 12075
rect 1105 11955 1145 11995
rect 1105 11875 1145 11915
rect 1105 11795 1145 11835
rect 1105 11715 1145 11755
rect 1105 11635 1145 11675
rect 1105 11555 1145 11595
rect 1105 11475 1145 11515
rect 1105 11395 1145 11435
rect 1105 11315 1145 11355
rect 1105 11235 1145 11275
rect 1105 11155 1145 11195
rect 1105 11075 1145 11115
rect 1105 10995 1145 11035
rect 1105 10915 1145 10955
rect 1105 10835 1145 10875
rect 1105 10755 1145 10795
rect 1105 10675 1145 10715
rect 1105 10595 1145 10635
rect 1105 10515 1145 10555
rect 1105 10435 1145 10475
rect 1105 10355 1145 10395
rect 1105 10275 1145 10315
rect 1220 12195 1260 12235
rect 1220 12115 1260 12155
rect 1220 12035 1260 12075
rect 1220 11955 1260 11995
rect 1220 11875 1260 11915
rect 1220 11795 1260 11835
rect 1220 11715 1260 11755
rect 1220 11635 1260 11675
rect 1220 11555 1260 11595
rect 1220 11475 1260 11515
rect 1220 11395 1260 11435
rect 1220 11315 1260 11355
rect 1220 11235 1260 11275
rect 1220 11155 1260 11195
rect 1220 11075 1260 11115
rect 1220 10995 1260 11035
rect 1220 10915 1260 10955
rect 1220 10835 1260 10875
rect 1220 10755 1260 10795
rect 1220 10675 1260 10715
rect 1220 10595 1260 10635
rect 1220 10515 1260 10555
rect 1220 10435 1260 10475
rect 1220 10355 1260 10395
rect 1220 10275 1260 10315
rect 1335 12195 1375 12235
rect 1335 12115 1375 12155
rect 1335 12035 1375 12075
rect 1335 11955 1375 11995
rect 1335 11875 1375 11915
rect 1335 11795 1375 11835
rect 1335 11715 1375 11755
rect 1335 11635 1375 11675
rect 1335 11555 1375 11595
rect 1335 11475 1375 11515
rect 1335 11395 1375 11435
rect 1335 11315 1375 11355
rect 1335 11235 1375 11275
rect 1335 11155 1375 11195
rect 1335 11075 1375 11115
rect 1335 10995 1375 11035
rect 1335 10915 1375 10955
rect 1335 10835 1375 10875
rect 1335 10755 1375 10795
rect 1335 10675 1375 10715
rect 1335 10595 1375 10635
rect 1335 10515 1375 10555
rect 1335 10435 1375 10475
rect 1335 10355 1375 10395
rect 1335 10275 1375 10315
rect 1450 12195 1490 12235
rect 1450 12115 1490 12155
rect 1450 12035 1490 12075
rect 1450 11955 1490 11995
rect 1450 11875 1490 11915
rect 1450 11795 1490 11835
rect 1450 11715 1490 11755
rect 1450 11635 1490 11675
rect 1450 11555 1490 11595
rect 1450 11475 1490 11515
rect 1450 11395 1490 11435
rect 1450 11315 1490 11355
rect 1450 11235 1490 11275
rect 1450 11155 1490 11195
rect 1450 11075 1490 11115
rect 1450 10995 1490 11035
rect 1450 10915 1490 10955
rect 1450 10835 1490 10875
rect 1450 10755 1490 10795
rect 1450 10675 1490 10715
rect 1450 10595 1490 10635
rect 1450 10515 1490 10555
rect 1450 10435 1490 10475
rect 1450 10355 1490 10395
rect 1450 10275 1490 10315
rect 1565 12195 1605 12235
rect 1565 12115 1605 12155
rect 1565 12035 1605 12075
rect 1565 11955 1605 11995
rect 1565 11875 1605 11915
rect 1565 11795 1605 11835
rect 1565 11715 1605 11755
rect 1565 11635 1605 11675
rect 1565 11555 1605 11595
rect 1565 11475 1605 11515
rect 1565 11395 1605 11435
rect 1565 11315 1605 11355
rect 1565 11235 1605 11275
rect 1565 11155 1605 11195
rect 1565 11075 1605 11115
rect 1565 10995 1605 11035
rect 1565 10915 1605 10955
rect 1565 10835 1605 10875
rect 1565 10755 1605 10795
rect 1565 10675 1605 10715
rect 1565 10595 1605 10635
rect 1565 10515 1605 10555
rect 1565 10435 1605 10475
rect 1565 10355 1605 10395
rect 1565 10275 1605 10315
rect 1680 12195 1720 12235
rect 1680 12115 1720 12155
rect 1680 12035 1720 12075
rect 1680 11955 1720 11995
rect 1680 11875 1720 11915
rect 1680 11795 1720 11835
rect 1680 11715 1720 11755
rect 1680 11635 1720 11675
rect 1680 11555 1720 11595
rect 1680 11475 1720 11515
rect 1680 11395 1720 11435
rect 1680 11315 1720 11355
rect 1680 11235 1720 11275
rect 1680 11155 1720 11195
rect 1680 11075 1720 11115
rect 1680 10995 1720 11035
rect 1680 10915 1720 10955
rect 1680 10835 1720 10875
rect 1680 10755 1720 10795
rect 1680 10675 1720 10715
rect 1680 10595 1720 10635
rect 1680 10515 1720 10555
rect 1680 10435 1720 10475
rect 1680 10355 1720 10395
rect 1680 10275 1720 10315
rect 1795 12195 1835 12235
rect 1795 12115 1835 12155
rect 1795 12035 1835 12075
rect 1795 11955 1835 11995
rect 1795 11875 1835 11915
rect 1795 11795 1835 11835
rect 1795 11715 1835 11755
rect 1795 11635 1835 11675
rect 1795 11555 1835 11595
rect 1795 11475 1835 11515
rect 1795 11395 1835 11435
rect 1795 11315 1835 11355
rect 1795 11235 1835 11275
rect 1795 11155 1835 11195
rect 1795 11075 1835 11115
rect 1795 10995 1835 11035
rect 1795 10915 1835 10955
rect 1795 10835 1835 10875
rect 1795 10755 1835 10795
rect 1795 10675 1835 10715
rect 1795 10595 1835 10635
rect 1795 10515 1835 10555
rect 1795 10435 1835 10475
rect 1795 10355 1835 10395
rect 1795 10275 1835 10315
rect 1910 12195 1950 12235
rect 1910 12115 1950 12155
rect 1910 12035 1950 12075
rect 1910 11955 1950 11995
rect 1910 11875 1950 11915
rect 1910 11795 1950 11835
rect 1910 11715 1950 11755
rect 1910 11635 1950 11675
rect 1910 11555 1950 11595
rect 1910 11475 1950 11515
rect 1910 11395 1950 11435
rect 1910 11315 1950 11355
rect 1910 11235 1950 11275
rect 1910 11155 1950 11195
rect 1910 11075 1950 11115
rect 1910 10995 1950 11035
rect 1910 10915 1950 10955
rect 1910 10835 1950 10875
rect 1910 10755 1950 10795
rect 1910 10675 1950 10715
rect 1910 10595 1950 10635
rect 1910 10515 1950 10555
rect 1910 10435 1950 10475
rect 1910 10355 1950 10395
rect 1910 10275 1950 10315
rect 2025 12195 2065 12235
rect 2025 12115 2065 12155
rect 2025 12035 2065 12075
rect 2025 11955 2065 11995
rect 2025 11875 2065 11915
rect 2025 11795 2065 11835
rect 2025 11715 2065 11755
rect 2025 11635 2065 11675
rect 2025 11555 2065 11595
rect 2025 11475 2065 11515
rect 2025 11395 2065 11435
rect 2025 11315 2065 11355
rect 2025 11235 2065 11275
rect 2025 11155 2065 11195
rect 2025 11075 2065 11115
rect 2025 10995 2065 11035
rect 2025 10915 2065 10955
rect 2025 10835 2065 10875
rect 2025 10755 2065 10795
rect 2025 10675 2065 10715
rect 2025 10595 2065 10635
rect 2025 10515 2065 10555
rect 2025 10435 2065 10475
rect 2025 10355 2065 10395
rect 2025 10275 2065 10315
rect 2140 12195 2180 12235
rect 2140 12115 2180 12155
rect 2140 12035 2180 12075
rect 2140 11955 2180 11995
rect 2140 11875 2180 11915
rect 2140 11795 2180 11835
rect 2140 11715 2180 11755
rect 2140 11635 2180 11675
rect 2140 11555 2180 11595
rect 2140 11475 2180 11515
rect 2140 11395 2180 11435
rect 2140 11315 2180 11355
rect 2140 11235 2180 11275
rect 2140 11155 2180 11195
rect 2140 11075 2180 11115
rect 2140 10995 2180 11035
rect 2140 10915 2180 10955
rect 2140 10835 2180 10875
rect 2140 10755 2180 10795
rect 2140 10675 2180 10715
rect 2140 10595 2180 10635
rect 2140 10515 2180 10555
rect 2140 10435 2180 10475
rect 2140 10355 2180 10395
rect 2140 10275 2180 10315
rect 2255 12195 2295 12235
rect 2255 12115 2295 12155
rect 2255 12035 2295 12075
rect 2255 11955 2295 11995
rect 2255 11875 2295 11915
rect 2255 11795 2295 11835
rect 2255 11715 2295 11755
rect 2255 11635 2295 11675
rect 2255 11555 2295 11595
rect 2255 11475 2295 11515
rect 2255 11395 2295 11435
rect 2255 11315 2295 11355
rect 2255 11235 2295 11275
rect 2255 11155 2295 11195
rect 2255 11075 2295 11115
rect 2255 10995 2295 11035
rect 2255 10915 2295 10955
rect 2255 10835 2295 10875
rect 2255 10755 2295 10795
rect 2255 10675 2295 10715
rect 2255 10595 2295 10635
rect 2255 10515 2295 10555
rect 2255 10435 2295 10475
rect 2255 10355 2295 10395
rect 2255 10275 2295 10315
rect 2370 12195 2410 12235
rect 2370 12115 2410 12155
rect 2370 12035 2410 12075
rect 2370 11955 2410 11995
rect 2370 11875 2410 11915
rect 2370 11795 2410 11835
rect 2370 11715 2410 11755
rect 2370 11635 2410 11675
rect 2370 11555 2410 11595
rect 2370 11475 2410 11515
rect 2370 11395 2410 11435
rect 2370 11315 2410 11355
rect 2370 11235 2410 11275
rect 2370 11155 2410 11195
rect 2370 11075 2410 11115
rect 2370 10995 2410 11035
rect 2370 10915 2410 10955
rect 2370 10835 2410 10875
rect 2370 10755 2410 10795
rect 2370 10675 2410 10715
rect 2370 10595 2410 10635
rect 2370 10515 2410 10555
rect 2370 10435 2410 10475
rect 2370 10355 2410 10395
rect 2370 10275 2410 10315
rect 2485 12195 2525 12235
rect 2485 12115 2525 12155
rect 2485 12035 2525 12075
rect 2485 11955 2525 11995
rect 2485 11875 2525 11915
rect 2485 11795 2525 11835
rect 2485 11715 2525 11755
rect 2485 11635 2525 11675
rect 2485 11555 2525 11595
rect 2485 11475 2525 11515
rect 2485 11395 2525 11435
rect 2485 11315 2525 11355
rect 2485 11235 2525 11275
rect 2485 11155 2525 11195
rect 2485 11075 2525 11115
rect 2485 10995 2525 11035
rect 2485 10915 2525 10955
rect 2485 10835 2525 10875
rect 2485 10755 2525 10795
rect 2485 10675 2525 10715
rect 2485 10595 2525 10635
rect 2485 10515 2525 10555
rect 2485 10435 2525 10475
rect 2485 10355 2525 10395
rect 2485 10275 2525 10315
rect 2685 12115 2725 12155
rect 2685 11955 2725 11995
rect 2685 11795 2725 11835
rect 2685 11635 2725 11675
rect 2685 11475 2725 11515
rect 2685 11315 2725 11355
rect 2685 11155 2725 11195
rect 2685 10915 2725 10955
rect 2685 10755 2725 10795
rect 2685 10595 2725 10635
rect 2685 10435 2725 10475
rect 2685 10275 2725 10315
rect -390 9990 -350 10030
rect -230 9990 -190 10030
rect -70 9990 -30 10030
rect 90 9990 130 10030
rect 250 9990 290 10030
rect 410 9990 450 10030
rect 570 9990 610 10030
rect 730 9990 770 10030
rect 1290 9990 1330 10030
rect 1450 9990 1490 10030
rect 1610 9990 1650 10030
rect 1770 9990 1810 10030
rect 1930 9990 1970 10030
rect 2090 9990 2130 10030
rect 2250 9990 2290 10030
rect 2410 9990 2450 10030
<< metal1 >>
rect -620 12475 880 12505
rect -620 12435 -390 12475
rect -350 12435 -230 12475
rect -190 12435 -70 12475
rect -30 12435 90 12475
rect 130 12435 250 12475
rect 290 12435 410 12475
rect 450 12435 570 12475
rect 610 12435 730 12475
rect 770 12435 880 12475
rect -620 12405 880 12435
rect 1265 12475 2755 12505
rect 1265 12435 1290 12475
rect 1330 12435 1450 12475
rect 1490 12435 1610 12475
rect 1650 12435 1770 12475
rect 1810 12435 1930 12475
rect 1970 12435 2090 12475
rect 2130 12435 2250 12475
rect 2290 12435 2410 12475
rect 2450 12435 2755 12475
rect 1265 12405 2755 12435
rect -1065 12340 3230 12370
rect -620 12235 -520 12285
rect -620 12195 -590 12235
rect -550 12195 -520 12235
rect -620 12075 -520 12195
rect -620 12035 -590 12075
rect -550 12035 -520 12075
rect -620 11915 -520 12035
rect -620 11875 -590 11915
rect -550 11875 -520 11915
rect -620 11755 -520 11875
rect -620 11715 -590 11755
rect -550 11715 -520 11755
rect -620 11595 -520 11715
rect -620 11555 -590 11595
rect -550 11555 -520 11595
rect -620 11435 -520 11555
rect -620 11395 -590 11435
rect -550 11395 -520 11435
rect -620 11275 -520 11395
rect -620 11235 -590 11275
rect -550 11235 -520 11275
rect -620 11115 -520 11235
rect -620 11075 -590 11115
rect -550 11075 -520 11115
rect -620 10955 -520 11075
rect -620 10915 -590 10955
rect -550 10915 -520 10955
rect -620 10795 -520 10915
rect -620 10755 -590 10795
rect -550 10755 -520 10795
rect -620 10635 -520 10755
rect -620 10595 -590 10635
rect -550 10595 -520 10635
rect -620 10475 -520 10595
rect -620 10435 -590 10475
rect -550 10435 -520 10475
rect -620 10315 -520 10435
rect -620 10275 -590 10315
rect -550 10275 -520 10315
rect -620 10230 -520 10275
rect -405 12255 -335 12340
rect -405 12235 -334 12255
rect -405 12195 -390 12235
rect -350 12195 -334 12235
rect -405 12155 -334 12195
rect -405 12115 -390 12155
rect -350 12115 -334 12155
rect -405 12075 -334 12115
rect -405 12035 -390 12075
rect -350 12035 -334 12075
rect -405 11995 -334 12035
rect -405 11955 -390 11995
rect -350 11955 -334 11995
rect -405 11915 -334 11955
rect -405 11875 -390 11915
rect -350 11875 -334 11915
rect -405 11835 -334 11875
rect -405 11795 -390 11835
rect -350 11795 -334 11835
rect -405 11755 -334 11795
rect -405 11715 -390 11755
rect -350 11715 -334 11755
rect -405 11675 -334 11715
rect -405 11635 -390 11675
rect -350 11635 -334 11675
rect -405 11595 -334 11635
rect -405 11555 -390 11595
rect -350 11555 -334 11595
rect -405 11515 -334 11555
rect -405 11475 -390 11515
rect -350 11475 -334 11515
rect -405 11435 -334 11475
rect -405 11395 -390 11435
rect -350 11395 -334 11435
rect -405 11355 -334 11395
rect -405 11315 -390 11355
rect -350 11315 -334 11355
rect -405 11275 -334 11315
rect -405 11235 -390 11275
rect -350 11235 -334 11275
rect -405 11195 -334 11235
rect -405 11155 -390 11195
rect -350 11155 -334 11195
rect -405 11115 -334 11155
rect -405 11075 -390 11115
rect -350 11075 -334 11115
rect -405 11035 -334 11075
rect -405 10995 -390 11035
rect -350 10995 -334 11035
rect -405 10955 -334 10995
rect -405 10915 -390 10955
rect -350 10915 -334 10955
rect -405 10875 -334 10915
rect -405 10835 -390 10875
rect -350 10835 -334 10875
rect -405 10795 -334 10835
rect -405 10755 -390 10795
rect -350 10755 -334 10795
rect -405 10715 -334 10755
rect -405 10675 -390 10715
rect -350 10675 -334 10715
rect -405 10635 -334 10675
rect -405 10595 -390 10635
rect -350 10595 -334 10635
rect -405 10555 -334 10595
rect -405 10515 -390 10555
rect -350 10515 -334 10555
rect -405 10475 -334 10515
rect -405 10435 -390 10475
rect -350 10435 -334 10475
rect -405 10395 -334 10435
rect -405 10355 -390 10395
rect -350 10355 -334 10395
rect -405 10315 -334 10355
rect -405 10275 -390 10315
rect -350 10275 -334 10315
rect -405 10260 -334 10275
rect -290 12235 -220 12255
rect -290 12195 -275 12235
rect -235 12195 -220 12235
rect -290 12155 -220 12195
rect -290 12115 -275 12155
rect -235 12115 -220 12155
rect -290 12075 -220 12115
rect -290 12035 -275 12075
rect -235 12035 -220 12075
rect -290 11995 -220 12035
rect -290 11955 -275 11995
rect -235 11955 -220 11995
rect -290 11915 -220 11955
rect -290 11875 -275 11915
rect -235 11875 -220 11915
rect -290 11835 -220 11875
rect -290 11795 -275 11835
rect -235 11795 -220 11835
rect -290 11755 -220 11795
rect -290 11715 -275 11755
rect -235 11715 -220 11755
rect -290 11675 -220 11715
rect -290 11635 -275 11675
rect -235 11635 -220 11675
rect -290 11595 -220 11635
rect -290 11555 -275 11595
rect -235 11555 -220 11595
rect -290 11515 -220 11555
rect -290 11475 -275 11515
rect -235 11475 -220 11515
rect -290 11435 -220 11475
rect -290 11395 -275 11435
rect -235 11395 -220 11435
rect -290 11355 -220 11395
rect -290 11315 -275 11355
rect -235 11315 -220 11355
rect -290 11275 -220 11315
rect -290 11235 -275 11275
rect -235 11235 -220 11275
rect -290 11195 -220 11235
rect -290 11155 -275 11195
rect -235 11155 -220 11195
rect -290 11115 -220 11155
rect -290 11075 -275 11115
rect -235 11075 -220 11115
rect -290 11035 -220 11075
rect -290 10995 -275 11035
rect -235 10995 -220 11035
rect -290 10955 -220 10995
rect -290 10915 -275 10955
rect -235 10915 -220 10955
rect -290 10875 -220 10915
rect -290 10835 -275 10875
rect -235 10835 -220 10875
rect -290 10795 -220 10835
rect -290 10755 -275 10795
rect -235 10755 -220 10795
rect -290 10715 -220 10755
rect -290 10675 -275 10715
rect -235 10675 -220 10715
rect -290 10635 -220 10675
rect -290 10595 -275 10635
rect -235 10595 -220 10635
rect -290 10555 -220 10595
rect -290 10515 -275 10555
rect -235 10515 -220 10555
rect -290 10475 -220 10515
rect -290 10435 -275 10475
rect -235 10435 -220 10475
rect -290 10395 -220 10435
rect -290 10355 -275 10395
rect -235 10355 -220 10395
rect -290 10315 -220 10355
rect -290 10275 -275 10315
rect -235 10275 -220 10315
rect -290 10150 -220 10275
rect -175 12235 -105 12340
rect -175 12195 -160 12235
rect -120 12195 -105 12235
rect -175 12155 -105 12195
rect -175 12115 -160 12155
rect -120 12115 -105 12155
rect -175 12075 -105 12115
rect -175 12035 -160 12075
rect -120 12035 -105 12075
rect -175 11995 -105 12035
rect -175 11955 -160 11995
rect -120 11955 -105 11995
rect -175 11915 -105 11955
rect -175 11875 -160 11915
rect -120 11875 -105 11915
rect -175 11835 -105 11875
rect -175 11795 -160 11835
rect -120 11795 -105 11835
rect -175 11755 -105 11795
rect -175 11715 -160 11755
rect -120 11715 -105 11755
rect -175 11675 -105 11715
rect -175 11635 -160 11675
rect -120 11635 -105 11675
rect -175 11595 -105 11635
rect -175 11555 -160 11595
rect -120 11555 -105 11595
rect -175 11515 -105 11555
rect -175 11475 -160 11515
rect -120 11475 -105 11515
rect -175 11435 -105 11475
rect -175 11395 -160 11435
rect -120 11395 -105 11435
rect -175 11355 -105 11395
rect -175 11315 -160 11355
rect -120 11315 -105 11355
rect -175 11275 -105 11315
rect -175 11235 -160 11275
rect -120 11235 -105 11275
rect -175 11195 -105 11235
rect -175 11155 -160 11195
rect -120 11155 -105 11195
rect -175 11115 -105 11155
rect -175 11075 -160 11115
rect -120 11075 -105 11115
rect -175 11035 -105 11075
rect -175 10995 -160 11035
rect -120 10995 -105 11035
rect -175 10955 -105 10995
rect -175 10915 -160 10955
rect -120 10915 -105 10955
rect -175 10875 -105 10915
rect -175 10835 -160 10875
rect -120 10835 -105 10875
rect -175 10795 -105 10835
rect -175 10755 -160 10795
rect -120 10755 -105 10795
rect -175 10715 -105 10755
rect -175 10675 -160 10715
rect -120 10675 -105 10715
rect -175 10635 -105 10675
rect -175 10595 -160 10635
rect -120 10595 -105 10635
rect -175 10555 -105 10595
rect -175 10515 -160 10555
rect -120 10515 -105 10555
rect -175 10475 -105 10515
rect -175 10435 -160 10475
rect -120 10435 -105 10475
rect -175 10395 -105 10435
rect -175 10355 -160 10395
rect -120 10355 -105 10395
rect -175 10315 -105 10355
rect -175 10275 -160 10315
rect -120 10275 -105 10315
rect -175 10260 -105 10275
rect -60 12235 10 12255
rect -60 12195 -45 12235
rect -5 12195 10 12235
rect -60 12155 10 12195
rect -60 12115 -45 12155
rect -5 12115 10 12155
rect -60 12075 10 12115
rect -60 12035 -45 12075
rect -5 12035 10 12075
rect -60 11995 10 12035
rect -60 11955 -45 11995
rect -5 11955 10 11995
rect -60 11915 10 11955
rect -60 11875 -45 11915
rect -5 11875 10 11915
rect -60 11835 10 11875
rect -60 11795 -45 11835
rect -5 11795 10 11835
rect -60 11755 10 11795
rect -60 11715 -45 11755
rect -5 11715 10 11755
rect -60 11675 10 11715
rect -60 11635 -45 11675
rect -5 11635 10 11675
rect -60 11595 10 11635
rect -60 11555 -45 11595
rect -5 11555 10 11595
rect -60 11515 10 11555
rect -60 11475 -45 11515
rect -5 11475 10 11515
rect -60 11435 10 11475
rect -60 11395 -45 11435
rect -5 11395 10 11435
rect -60 11355 10 11395
rect -60 11315 -45 11355
rect -5 11315 10 11355
rect -60 11275 10 11315
rect -60 11235 -45 11275
rect -5 11235 10 11275
rect -60 11195 10 11235
rect -60 11155 -45 11195
rect -5 11155 10 11195
rect -60 11115 10 11155
rect -60 11075 -45 11115
rect -5 11075 10 11115
rect -60 11035 10 11075
rect -60 10995 -45 11035
rect -5 10995 10 11035
rect -60 10955 10 10995
rect -60 10915 -45 10955
rect -5 10915 10 10955
rect -60 10875 10 10915
rect -60 10835 -45 10875
rect -5 10835 10 10875
rect -60 10795 10 10835
rect -60 10755 -45 10795
rect -5 10755 10 10795
rect -60 10715 10 10755
rect -60 10675 -45 10715
rect -5 10675 10 10715
rect -60 10635 10 10675
rect -60 10595 -45 10635
rect -5 10595 10 10635
rect -60 10555 10 10595
rect -60 10515 -45 10555
rect -5 10515 10 10555
rect -60 10475 10 10515
rect -60 10435 -45 10475
rect -5 10435 10 10475
rect -60 10395 10 10435
rect -60 10355 -45 10395
rect -5 10355 10 10395
rect -60 10315 10 10355
rect -60 10275 -45 10315
rect -5 10275 10 10315
rect -60 10150 10 10275
rect 55 12235 125 12340
rect 55 12195 70 12235
rect 110 12195 125 12235
rect 55 12155 125 12195
rect 55 12115 70 12155
rect 110 12115 125 12155
rect 55 12075 125 12115
rect 55 12035 70 12075
rect 110 12035 125 12075
rect 55 11995 125 12035
rect 55 11955 70 11995
rect 110 11955 125 11995
rect 55 11915 125 11955
rect 55 11875 70 11915
rect 110 11875 125 11915
rect 55 11835 125 11875
rect 55 11795 70 11835
rect 110 11795 125 11835
rect 55 11755 125 11795
rect 55 11715 70 11755
rect 110 11715 125 11755
rect 55 11675 125 11715
rect 55 11635 70 11675
rect 110 11635 125 11675
rect 55 11595 125 11635
rect 55 11555 70 11595
rect 110 11555 125 11595
rect 55 11515 125 11555
rect 55 11475 70 11515
rect 110 11475 125 11515
rect 55 11435 125 11475
rect 55 11395 70 11435
rect 110 11395 125 11435
rect 55 11355 125 11395
rect 55 11315 70 11355
rect 110 11315 125 11355
rect 55 11275 125 11315
rect 55 11235 70 11275
rect 110 11235 125 11275
rect 55 11195 125 11235
rect 55 11155 70 11195
rect 110 11155 125 11195
rect 55 11115 125 11155
rect 55 11075 70 11115
rect 110 11075 125 11115
rect 55 11035 125 11075
rect 55 10995 70 11035
rect 110 10995 125 11035
rect 55 10955 125 10995
rect 55 10915 70 10955
rect 110 10915 125 10955
rect 55 10875 125 10915
rect 55 10835 70 10875
rect 110 10835 125 10875
rect 55 10795 125 10835
rect 55 10755 70 10795
rect 110 10755 125 10795
rect 55 10715 125 10755
rect 55 10675 70 10715
rect 110 10675 125 10715
rect 55 10635 125 10675
rect 55 10595 70 10635
rect 110 10595 125 10635
rect 55 10555 125 10595
rect 55 10515 70 10555
rect 110 10515 125 10555
rect 55 10475 125 10515
rect 55 10435 70 10475
rect 110 10435 125 10475
rect 55 10395 125 10435
rect 55 10355 70 10395
rect 110 10355 125 10395
rect 55 10315 125 10355
rect 55 10275 70 10315
rect 110 10275 125 10315
rect 55 10260 125 10275
rect 170 12235 240 12255
rect 170 12195 185 12235
rect 225 12195 240 12235
rect 170 12155 240 12195
rect 170 12115 185 12155
rect 225 12115 240 12155
rect 170 12075 240 12115
rect 170 12035 185 12075
rect 225 12035 240 12075
rect 170 11995 240 12035
rect 170 11955 185 11995
rect 225 11955 240 11995
rect 170 11915 240 11955
rect 170 11875 185 11915
rect 225 11875 240 11915
rect 170 11835 240 11875
rect 170 11795 185 11835
rect 225 11795 240 11835
rect 170 11755 240 11795
rect 170 11715 185 11755
rect 225 11715 240 11755
rect 170 11675 240 11715
rect 170 11635 185 11675
rect 225 11635 240 11675
rect 170 11595 240 11635
rect 170 11555 185 11595
rect 225 11555 240 11595
rect 170 11515 240 11555
rect 170 11475 185 11515
rect 225 11475 240 11515
rect 170 11435 240 11475
rect 170 11395 185 11435
rect 225 11395 240 11435
rect 170 11355 240 11395
rect 170 11315 185 11355
rect 225 11315 240 11355
rect 170 11275 240 11315
rect 170 11235 185 11275
rect 225 11235 240 11275
rect 170 11195 240 11235
rect 170 11155 185 11195
rect 225 11155 240 11195
rect 170 11115 240 11155
rect 170 11075 185 11115
rect 225 11075 240 11115
rect 170 11035 240 11075
rect 170 10995 185 11035
rect 225 10995 240 11035
rect 170 10955 240 10995
rect 170 10915 185 10955
rect 225 10915 240 10955
rect 170 10875 240 10915
rect 170 10835 185 10875
rect 225 10835 240 10875
rect 170 10795 240 10835
rect 170 10755 185 10795
rect 225 10755 240 10795
rect 170 10715 240 10755
rect 170 10675 185 10715
rect 225 10675 240 10715
rect 170 10635 240 10675
rect 170 10595 185 10635
rect 225 10595 240 10635
rect 170 10555 240 10595
rect 170 10515 185 10555
rect 225 10515 240 10555
rect 170 10475 240 10515
rect 170 10435 185 10475
rect 225 10435 240 10475
rect 170 10395 240 10435
rect 170 10355 185 10395
rect 225 10355 240 10395
rect 170 10315 240 10355
rect 170 10275 185 10315
rect 225 10275 240 10315
rect 170 10150 240 10275
rect 285 12235 355 12340
rect 285 12195 300 12235
rect 340 12195 355 12235
rect 285 12155 355 12195
rect 285 12115 300 12155
rect 340 12115 355 12155
rect 285 12075 355 12115
rect 285 12035 300 12075
rect 340 12035 355 12075
rect 285 11995 355 12035
rect 285 11955 300 11995
rect 340 11955 355 11995
rect 285 11915 355 11955
rect 285 11875 300 11915
rect 340 11875 355 11915
rect 285 11835 355 11875
rect 285 11795 300 11835
rect 340 11795 355 11835
rect 285 11755 355 11795
rect 285 11715 300 11755
rect 340 11715 355 11755
rect 285 11675 355 11715
rect 285 11635 300 11675
rect 340 11635 355 11675
rect 285 11595 355 11635
rect 285 11555 300 11595
rect 340 11555 355 11595
rect 285 11515 355 11555
rect 285 11475 300 11515
rect 340 11475 355 11515
rect 285 11435 355 11475
rect 285 11395 300 11435
rect 340 11395 355 11435
rect 285 11355 355 11395
rect 285 11315 300 11355
rect 340 11315 355 11355
rect 285 11275 355 11315
rect 285 11235 300 11275
rect 340 11235 355 11275
rect 285 11195 355 11235
rect 285 11155 300 11195
rect 340 11155 355 11195
rect 285 11115 355 11155
rect 285 11075 300 11115
rect 340 11075 355 11115
rect 285 11035 355 11075
rect 285 10995 300 11035
rect 340 10995 355 11035
rect 285 10955 355 10995
rect 285 10915 300 10955
rect 340 10915 355 10955
rect 285 10875 355 10915
rect 285 10835 300 10875
rect 340 10835 355 10875
rect 285 10795 355 10835
rect 285 10755 300 10795
rect 340 10755 355 10795
rect 285 10715 355 10755
rect 285 10675 300 10715
rect 340 10675 355 10715
rect 285 10635 355 10675
rect 285 10595 300 10635
rect 340 10595 355 10635
rect 285 10555 355 10595
rect 285 10515 300 10555
rect 340 10515 355 10555
rect 285 10475 355 10515
rect 285 10435 300 10475
rect 340 10435 355 10475
rect 285 10395 355 10435
rect 285 10355 300 10395
rect 340 10355 355 10395
rect 285 10315 355 10355
rect 285 10275 300 10315
rect 340 10275 355 10315
rect 285 10260 355 10275
rect 400 12235 470 12255
rect 400 12195 415 12235
rect 455 12195 470 12235
rect 400 12155 470 12195
rect 400 12115 415 12155
rect 455 12115 470 12155
rect 400 12075 470 12115
rect 400 12035 415 12075
rect 455 12035 470 12075
rect 400 11995 470 12035
rect 400 11955 415 11995
rect 455 11955 470 11995
rect 400 11915 470 11955
rect 400 11875 415 11915
rect 455 11875 470 11915
rect 400 11835 470 11875
rect 400 11795 415 11835
rect 455 11795 470 11835
rect 400 11755 470 11795
rect 400 11715 415 11755
rect 455 11715 470 11755
rect 400 11675 470 11715
rect 400 11635 415 11675
rect 455 11635 470 11675
rect 400 11595 470 11635
rect 400 11555 415 11595
rect 455 11555 470 11595
rect 400 11515 470 11555
rect 400 11475 415 11515
rect 455 11475 470 11515
rect 400 11435 470 11475
rect 400 11395 415 11435
rect 455 11395 470 11435
rect 400 11355 470 11395
rect 400 11315 415 11355
rect 455 11315 470 11355
rect 400 11275 470 11315
rect 400 11235 415 11275
rect 455 11235 470 11275
rect 400 11195 470 11235
rect 400 11155 415 11195
rect 455 11155 470 11195
rect 400 11115 470 11155
rect 400 11075 415 11115
rect 455 11075 470 11115
rect 400 11035 470 11075
rect 400 10995 415 11035
rect 455 10995 470 11035
rect 400 10955 470 10995
rect 400 10915 415 10955
rect 455 10915 470 10955
rect 400 10875 470 10915
rect 400 10835 415 10875
rect 455 10835 470 10875
rect 400 10795 470 10835
rect 400 10755 415 10795
rect 455 10755 470 10795
rect 400 10715 470 10755
rect 400 10675 415 10715
rect 455 10675 470 10715
rect 400 10635 470 10675
rect 400 10595 415 10635
rect 455 10595 470 10635
rect 400 10555 470 10595
rect 400 10515 415 10555
rect 455 10515 470 10555
rect 400 10475 470 10515
rect 400 10435 415 10475
rect 455 10435 470 10475
rect 400 10395 470 10435
rect 400 10355 415 10395
rect 455 10355 470 10395
rect 400 10315 470 10355
rect 400 10275 415 10315
rect 455 10275 470 10315
rect 400 10150 470 10275
rect 515 12235 585 12340
rect 515 12195 530 12235
rect 570 12195 585 12235
rect 515 12155 585 12195
rect 515 12115 530 12155
rect 570 12115 585 12155
rect 515 12075 585 12115
rect 515 12035 530 12075
rect 570 12035 585 12075
rect 515 11995 585 12035
rect 515 11955 530 11995
rect 570 11955 585 11995
rect 515 11915 585 11955
rect 515 11875 530 11915
rect 570 11875 585 11915
rect 515 11835 585 11875
rect 515 11795 530 11835
rect 570 11795 585 11835
rect 515 11755 585 11795
rect 515 11715 530 11755
rect 570 11715 585 11755
rect 515 11675 585 11715
rect 515 11635 530 11675
rect 570 11635 585 11675
rect 515 11595 585 11635
rect 515 11555 530 11595
rect 570 11555 585 11595
rect 515 11515 585 11555
rect 515 11475 530 11515
rect 570 11475 585 11515
rect 515 11435 585 11475
rect 515 11395 530 11435
rect 570 11395 585 11435
rect 515 11355 585 11395
rect 515 11315 530 11355
rect 570 11315 585 11355
rect 515 11275 585 11315
rect 515 11235 530 11275
rect 570 11235 585 11275
rect 515 11195 585 11235
rect 515 11155 530 11195
rect 570 11155 585 11195
rect 515 11115 585 11155
rect 515 11075 530 11115
rect 570 11075 585 11115
rect 515 11035 585 11075
rect 515 10995 530 11035
rect 570 10995 585 11035
rect 515 10955 585 10995
rect 515 10915 530 10955
rect 570 10915 585 10955
rect 515 10875 585 10915
rect 515 10835 530 10875
rect 570 10835 585 10875
rect 515 10795 585 10835
rect 515 10755 530 10795
rect 570 10755 585 10795
rect 515 10715 585 10755
rect 515 10675 530 10715
rect 570 10675 585 10715
rect 515 10635 585 10675
rect 515 10595 530 10635
rect 570 10595 585 10635
rect 515 10555 585 10595
rect 515 10515 530 10555
rect 570 10515 585 10555
rect 515 10475 585 10515
rect 515 10435 530 10475
rect 570 10435 585 10475
rect 515 10395 585 10435
rect 515 10355 530 10395
rect 570 10355 585 10395
rect 515 10315 585 10355
rect 515 10275 530 10315
rect 570 10275 585 10315
rect 515 10260 585 10275
rect 630 12235 700 12255
rect 630 12195 645 12235
rect 685 12195 700 12235
rect 630 12155 700 12195
rect 630 12115 645 12155
rect 685 12115 700 12155
rect 630 12075 700 12115
rect 630 12035 645 12075
rect 685 12035 700 12075
rect 630 11995 700 12035
rect 630 11955 645 11995
rect 685 11955 700 11995
rect 630 11915 700 11955
rect 630 11875 645 11915
rect 685 11875 700 11915
rect 630 11835 700 11875
rect 630 11795 645 11835
rect 685 11795 700 11835
rect 630 11755 700 11795
rect 630 11715 645 11755
rect 685 11715 700 11755
rect 630 11675 700 11715
rect 630 11635 645 11675
rect 685 11635 700 11675
rect 630 11595 700 11635
rect 630 11555 645 11595
rect 685 11555 700 11595
rect 630 11515 700 11555
rect 630 11475 645 11515
rect 685 11475 700 11515
rect 630 11435 700 11475
rect 630 11395 645 11435
rect 685 11395 700 11435
rect 630 11355 700 11395
rect 630 11315 645 11355
rect 685 11315 700 11355
rect 630 11275 700 11315
rect 630 11235 645 11275
rect 685 11235 700 11275
rect 630 11195 700 11235
rect 630 11155 645 11195
rect 685 11155 700 11195
rect 630 11115 700 11155
rect 630 11075 645 11115
rect 685 11075 700 11115
rect 630 11035 700 11075
rect 630 10995 645 11035
rect 685 10995 700 11035
rect 630 10955 700 10995
rect 630 10915 645 10955
rect 685 10915 700 10955
rect 630 10875 700 10915
rect 630 10835 645 10875
rect 685 10835 700 10875
rect 630 10795 700 10835
rect 630 10755 645 10795
rect 685 10755 700 10795
rect 630 10715 700 10755
rect 630 10675 645 10715
rect 685 10675 700 10715
rect 630 10635 700 10675
rect 630 10595 645 10635
rect 685 10595 700 10635
rect 630 10555 700 10595
rect 630 10515 645 10555
rect 685 10515 700 10555
rect 630 10475 700 10515
rect 630 10435 645 10475
rect 685 10435 700 10475
rect 630 10395 700 10435
rect 630 10355 645 10395
rect 685 10355 700 10395
rect 630 10315 700 10355
rect 630 10275 645 10315
rect 685 10275 700 10315
rect 630 10150 700 10275
rect 745 12235 815 12340
rect 745 12195 760 12235
rect 800 12195 815 12235
rect 745 12155 815 12195
rect 745 12115 760 12155
rect 800 12115 815 12155
rect 745 12075 815 12115
rect 745 12035 760 12075
rect 800 12035 815 12075
rect 745 11995 815 12035
rect 745 11955 760 11995
rect 800 11955 815 11995
rect 745 11915 815 11955
rect 745 11875 760 11915
rect 800 11875 815 11915
rect 745 11835 815 11875
rect 745 11795 760 11835
rect 800 11795 815 11835
rect 745 11755 815 11795
rect 745 11715 760 11755
rect 800 11715 815 11755
rect 745 11675 815 11715
rect 745 11635 760 11675
rect 800 11635 815 11675
rect 745 11595 815 11635
rect 745 11555 760 11595
rect 800 11555 815 11595
rect 745 11515 815 11555
rect 745 11475 760 11515
rect 800 11475 815 11515
rect 745 11435 815 11475
rect 745 11395 760 11435
rect 800 11395 815 11435
rect 745 11355 815 11395
rect 745 11315 760 11355
rect 800 11315 815 11355
rect 745 11275 815 11315
rect 745 11235 760 11275
rect 800 11235 815 11275
rect 745 11195 815 11235
rect 745 11155 760 11195
rect 800 11155 815 11195
rect 745 11115 815 11155
rect 745 11075 760 11115
rect 800 11075 815 11115
rect 745 11035 815 11075
rect 745 10995 760 11035
rect 800 10995 815 11035
rect 745 10955 815 10995
rect 745 10915 760 10955
rect 800 10915 815 10955
rect 745 10875 815 10915
rect 745 10835 760 10875
rect 800 10835 815 10875
rect 745 10795 815 10835
rect 745 10755 760 10795
rect 800 10755 815 10795
rect 745 10715 815 10755
rect 745 10675 760 10715
rect 800 10675 815 10715
rect 745 10635 815 10675
rect 745 10595 760 10635
rect 800 10595 815 10635
rect 745 10555 815 10595
rect 745 10515 760 10555
rect 800 10515 815 10555
rect 745 10475 815 10515
rect 745 10435 760 10475
rect 800 10435 815 10475
rect 745 10395 815 10435
rect 745 10355 760 10395
rect 800 10355 815 10395
rect 745 10315 815 10355
rect 745 10275 760 10315
rect 800 10275 815 10315
rect 745 10260 815 10275
rect 860 12235 930 12255
rect 860 12195 875 12235
rect 915 12195 930 12235
rect 860 12155 930 12195
rect 860 12115 875 12155
rect 915 12115 930 12155
rect 860 12075 930 12115
rect 860 12035 875 12075
rect 915 12035 930 12075
rect 860 11995 930 12035
rect 860 11955 875 11995
rect 915 11955 930 11995
rect 860 11915 930 11955
rect 860 11875 875 11915
rect 915 11875 930 11915
rect 860 11835 930 11875
rect 860 11795 875 11835
rect 915 11795 930 11835
rect 860 11755 930 11795
rect 860 11715 875 11755
rect 915 11715 930 11755
rect 860 11675 930 11715
rect 860 11635 875 11675
rect 915 11635 930 11675
rect 860 11595 930 11635
rect 860 11555 875 11595
rect 915 11555 930 11595
rect 860 11515 930 11555
rect 860 11475 875 11515
rect 915 11475 930 11515
rect 860 11435 930 11475
rect 860 11395 875 11435
rect 915 11395 930 11435
rect 860 11355 930 11395
rect 860 11315 875 11355
rect 915 11315 930 11355
rect 860 11275 930 11315
rect 860 11235 875 11275
rect 915 11235 930 11275
rect 860 11195 930 11235
rect 860 11155 875 11195
rect 915 11155 930 11195
rect 860 11115 930 11155
rect 860 11075 875 11115
rect 915 11075 930 11115
rect 860 11035 930 11075
rect 860 10995 875 11035
rect 915 10995 930 11035
rect 860 10955 930 10995
rect 860 10915 875 10955
rect 915 10915 930 10955
rect 860 10875 930 10915
rect 860 10835 875 10875
rect 915 10835 930 10875
rect 860 10795 930 10835
rect 860 10755 875 10795
rect 915 10755 930 10795
rect 860 10715 930 10755
rect 860 10675 875 10715
rect 915 10675 930 10715
rect 860 10635 930 10675
rect 860 10595 875 10635
rect 915 10595 930 10635
rect 860 10555 930 10595
rect 860 10515 875 10555
rect 915 10515 930 10555
rect 860 10475 930 10515
rect 860 10435 875 10475
rect 915 10435 930 10475
rect 860 10395 930 10435
rect 860 10355 875 10395
rect 915 10355 930 10395
rect 860 10315 930 10355
rect 860 10275 875 10315
rect 915 10275 930 10315
rect 860 10150 930 10275
rect 975 12235 1045 12340
rect 975 12195 990 12235
rect 1030 12195 1045 12235
rect 975 12155 1045 12195
rect 975 12115 990 12155
rect 1030 12115 1045 12155
rect 975 12075 1045 12115
rect 975 12035 990 12075
rect 1030 12035 1045 12075
rect 975 11995 1045 12035
rect 975 11955 990 11995
rect 1030 11955 1045 11995
rect 975 11915 1045 11955
rect 975 11875 990 11915
rect 1030 11875 1045 11915
rect 975 11835 1045 11875
rect 975 11795 990 11835
rect 1030 11795 1045 11835
rect 975 11755 1045 11795
rect 975 11715 990 11755
rect 1030 11715 1045 11755
rect 975 11675 1045 11715
rect 975 11635 990 11675
rect 1030 11635 1045 11675
rect 975 11595 1045 11635
rect 975 11555 990 11595
rect 1030 11555 1045 11595
rect 975 11515 1045 11555
rect 975 11475 990 11515
rect 1030 11475 1045 11515
rect 975 11435 1045 11475
rect 975 11395 990 11435
rect 1030 11395 1045 11435
rect 975 11355 1045 11395
rect 975 11315 990 11355
rect 1030 11315 1045 11355
rect 975 11275 1045 11315
rect 975 11235 990 11275
rect 1030 11235 1045 11275
rect 975 11195 1045 11235
rect 975 11155 990 11195
rect 1030 11155 1045 11195
rect 975 11115 1045 11155
rect 975 11075 990 11115
rect 1030 11075 1045 11115
rect 975 11035 1045 11075
rect 975 10995 990 11035
rect 1030 10995 1045 11035
rect 975 10955 1045 10995
rect 975 10915 990 10955
rect 1030 10915 1045 10955
rect 975 10875 1045 10915
rect 975 10835 990 10875
rect 1030 10835 1045 10875
rect 975 10795 1045 10835
rect 975 10755 990 10795
rect 1030 10755 1045 10795
rect 975 10715 1045 10755
rect 975 10675 990 10715
rect 1030 10675 1045 10715
rect 975 10635 1045 10675
rect 975 10595 990 10635
rect 1030 10595 1045 10635
rect 975 10555 1045 10595
rect 975 10515 990 10555
rect 1030 10515 1045 10555
rect 975 10475 1045 10515
rect 975 10435 990 10475
rect 1030 10435 1045 10475
rect 975 10395 1045 10435
rect 975 10355 990 10395
rect 1030 10355 1045 10395
rect 975 10315 1045 10355
rect 975 10275 990 10315
rect 1030 10275 1045 10315
rect 975 10260 1045 10275
rect 1090 12235 1160 12255
rect 1090 12195 1105 12235
rect 1145 12195 1160 12235
rect 1090 12155 1160 12195
rect 1090 12115 1105 12155
rect 1145 12115 1160 12155
rect 1090 12075 1160 12115
rect 1090 12035 1105 12075
rect 1145 12035 1160 12075
rect 1090 11995 1160 12035
rect 1090 11955 1105 11995
rect 1145 11955 1160 11995
rect 1090 11915 1160 11955
rect 1090 11875 1105 11915
rect 1145 11875 1160 11915
rect 1090 11835 1160 11875
rect 1090 11795 1105 11835
rect 1145 11795 1160 11835
rect 1090 11755 1160 11795
rect 1090 11715 1105 11755
rect 1145 11715 1160 11755
rect 1090 11675 1160 11715
rect 1090 11635 1105 11675
rect 1145 11635 1160 11675
rect 1090 11595 1160 11635
rect 1090 11555 1105 11595
rect 1145 11555 1160 11595
rect 1090 11515 1160 11555
rect 1090 11475 1105 11515
rect 1145 11475 1160 11515
rect 1090 11435 1160 11475
rect 1090 11395 1105 11435
rect 1145 11395 1160 11435
rect 1090 11355 1160 11395
rect 1090 11315 1105 11355
rect 1145 11315 1160 11355
rect 1090 11275 1160 11315
rect 1090 11235 1105 11275
rect 1145 11235 1160 11275
rect 1090 11195 1160 11235
rect 1090 11155 1105 11195
rect 1145 11155 1160 11195
rect 1090 11115 1160 11155
rect 1090 11075 1105 11115
rect 1145 11075 1160 11115
rect 1090 11035 1160 11075
rect 1090 10995 1105 11035
rect 1145 10995 1160 11035
rect 1090 10955 1160 10995
rect 1090 10915 1105 10955
rect 1145 10915 1160 10955
rect 1090 10875 1160 10915
rect 1090 10835 1105 10875
rect 1145 10835 1160 10875
rect 1090 10795 1160 10835
rect 1090 10755 1105 10795
rect 1145 10755 1160 10795
rect 1090 10715 1160 10755
rect 1090 10675 1105 10715
rect 1145 10675 1160 10715
rect 1090 10635 1160 10675
rect 1090 10595 1105 10635
rect 1145 10595 1160 10635
rect 1090 10555 1160 10595
rect 1090 10515 1105 10555
rect 1145 10515 1160 10555
rect 1090 10475 1160 10515
rect 1090 10435 1105 10475
rect 1145 10435 1160 10475
rect 1090 10395 1160 10435
rect 1090 10355 1105 10395
rect 1145 10355 1160 10395
rect 1090 10315 1160 10355
rect 1090 10275 1105 10315
rect 1145 10275 1160 10315
rect 1090 10150 1160 10275
rect 1205 12235 1275 12340
rect 1205 12195 1220 12235
rect 1260 12195 1275 12235
rect 1205 12155 1275 12195
rect 1205 12115 1220 12155
rect 1260 12115 1275 12155
rect 1205 12075 1275 12115
rect 1205 12035 1220 12075
rect 1260 12035 1275 12075
rect 1205 11995 1275 12035
rect 1205 11955 1220 11995
rect 1260 11955 1275 11995
rect 1205 11915 1275 11955
rect 1205 11875 1220 11915
rect 1260 11875 1275 11915
rect 1205 11835 1275 11875
rect 1205 11795 1220 11835
rect 1260 11795 1275 11835
rect 1205 11755 1275 11795
rect 1205 11715 1220 11755
rect 1260 11715 1275 11755
rect 1205 11675 1275 11715
rect 1205 11635 1220 11675
rect 1260 11635 1275 11675
rect 1205 11595 1275 11635
rect 1205 11555 1220 11595
rect 1260 11555 1275 11595
rect 1205 11515 1275 11555
rect 1205 11475 1220 11515
rect 1260 11475 1275 11515
rect 1205 11435 1275 11475
rect 1205 11395 1220 11435
rect 1260 11395 1275 11435
rect 1205 11355 1275 11395
rect 1205 11315 1220 11355
rect 1260 11315 1275 11355
rect 1205 11275 1275 11315
rect 1205 11235 1220 11275
rect 1260 11235 1275 11275
rect 1205 11195 1275 11235
rect 1205 11155 1220 11195
rect 1260 11155 1275 11195
rect 1205 11115 1275 11155
rect 1205 11075 1220 11115
rect 1260 11075 1275 11115
rect 1205 11035 1275 11075
rect 1205 10995 1220 11035
rect 1260 10995 1275 11035
rect 1205 10955 1275 10995
rect 1205 10915 1220 10955
rect 1260 10915 1275 10955
rect 1205 10875 1275 10915
rect 1205 10835 1220 10875
rect 1260 10835 1275 10875
rect 1205 10795 1275 10835
rect 1205 10755 1220 10795
rect 1260 10755 1275 10795
rect 1205 10715 1275 10755
rect 1205 10675 1220 10715
rect 1260 10675 1275 10715
rect 1205 10635 1275 10675
rect 1205 10595 1220 10635
rect 1260 10595 1275 10635
rect 1205 10555 1275 10595
rect 1205 10515 1220 10555
rect 1260 10515 1275 10555
rect 1205 10475 1275 10515
rect 1205 10435 1220 10475
rect 1260 10435 1275 10475
rect 1205 10395 1275 10435
rect 1205 10355 1220 10395
rect 1260 10355 1275 10395
rect 1205 10315 1275 10355
rect 1205 10275 1220 10315
rect 1260 10275 1275 10315
rect 1205 10260 1275 10275
rect 1320 12235 1390 12255
rect 1320 12195 1335 12235
rect 1375 12195 1390 12235
rect 1320 12155 1390 12195
rect 1320 12115 1335 12155
rect 1375 12115 1390 12155
rect 1320 12075 1390 12115
rect 1320 12035 1335 12075
rect 1375 12035 1390 12075
rect 1320 11995 1390 12035
rect 1320 11955 1335 11995
rect 1375 11955 1390 11995
rect 1320 11915 1390 11955
rect 1320 11875 1335 11915
rect 1375 11875 1390 11915
rect 1320 11835 1390 11875
rect 1320 11795 1335 11835
rect 1375 11795 1390 11835
rect 1320 11755 1390 11795
rect 1320 11715 1335 11755
rect 1375 11715 1390 11755
rect 1320 11675 1390 11715
rect 1320 11635 1335 11675
rect 1375 11635 1390 11675
rect 1320 11595 1390 11635
rect 1320 11555 1335 11595
rect 1375 11555 1390 11595
rect 1320 11515 1390 11555
rect 1320 11475 1335 11515
rect 1375 11475 1390 11515
rect 1320 11435 1390 11475
rect 1320 11395 1335 11435
rect 1375 11395 1390 11435
rect 1320 11355 1390 11395
rect 1320 11315 1335 11355
rect 1375 11315 1390 11355
rect 1320 11275 1390 11315
rect 1320 11235 1335 11275
rect 1375 11235 1390 11275
rect 1320 11195 1390 11235
rect 1320 11155 1335 11195
rect 1375 11155 1390 11195
rect 1320 11115 1390 11155
rect 1320 11075 1335 11115
rect 1375 11075 1390 11115
rect 1320 11035 1390 11075
rect 1320 10995 1335 11035
rect 1375 10995 1390 11035
rect 1320 10955 1390 10995
rect 1320 10915 1335 10955
rect 1375 10915 1390 10955
rect 1320 10875 1390 10915
rect 1320 10835 1335 10875
rect 1375 10835 1390 10875
rect 1320 10795 1390 10835
rect 1320 10755 1335 10795
rect 1375 10755 1390 10795
rect 1320 10715 1390 10755
rect 1320 10675 1335 10715
rect 1375 10675 1390 10715
rect 1320 10635 1390 10675
rect 1320 10595 1335 10635
rect 1375 10595 1390 10635
rect 1320 10555 1390 10595
rect 1320 10515 1335 10555
rect 1375 10515 1390 10555
rect 1320 10475 1390 10515
rect 1320 10435 1335 10475
rect 1375 10435 1390 10475
rect 1320 10395 1390 10435
rect 1320 10355 1335 10395
rect 1375 10355 1390 10395
rect 1320 10315 1390 10355
rect 1320 10275 1335 10315
rect 1375 10275 1390 10315
rect 1320 10150 1390 10275
rect 1435 12235 1505 12340
rect 1435 12195 1450 12235
rect 1490 12195 1505 12235
rect 1435 12155 1505 12195
rect 1435 12115 1450 12155
rect 1490 12115 1505 12155
rect 1435 12075 1505 12115
rect 1435 12035 1450 12075
rect 1490 12035 1505 12075
rect 1435 11995 1505 12035
rect 1435 11955 1450 11995
rect 1490 11955 1505 11995
rect 1435 11915 1505 11955
rect 1435 11875 1450 11915
rect 1490 11875 1505 11915
rect 1435 11835 1505 11875
rect 1435 11795 1450 11835
rect 1490 11795 1505 11835
rect 1435 11755 1505 11795
rect 1435 11715 1450 11755
rect 1490 11715 1505 11755
rect 1435 11675 1505 11715
rect 1435 11635 1450 11675
rect 1490 11635 1505 11675
rect 1435 11595 1505 11635
rect 1435 11555 1450 11595
rect 1490 11555 1505 11595
rect 1435 11515 1505 11555
rect 1435 11475 1450 11515
rect 1490 11475 1505 11515
rect 1435 11435 1505 11475
rect 1435 11395 1450 11435
rect 1490 11395 1505 11435
rect 1435 11355 1505 11395
rect 1435 11315 1450 11355
rect 1490 11315 1505 11355
rect 1435 11275 1505 11315
rect 1435 11235 1450 11275
rect 1490 11235 1505 11275
rect 1435 11195 1505 11235
rect 1435 11155 1450 11195
rect 1490 11155 1505 11195
rect 1435 11115 1505 11155
rect 1435 11075 1450 11115
rect 1490 11075 1505 11115
rect 1435 11035 1505 11075
rect 1435 10995 1450 11035
rect 1490 10995 1505 11035
rect 1435 10955 1505 10995
rect 1435 10915 1450 10955
rect 1490 10915 1505 10955
rect 1435 10875 1505 10915
rect 1435 10835 1450 10875
rect 1490 10835 1505 10875
rect 1435 10795 1505 10835
rect 1435 10755 1450 10795
rect 1490 10755 1505 10795
rect 1435 10715 1505 10755
rect 1435 10675 1450 10715
rect 1490 10675 1505 10715
rect 1435 10635 1505 10675
rect 1435 10595 1450 10635
rect 1490 10595 1505 10635
rect 1435 10555 1505 10595
rect 1435 10515 1450 10555
rect 1490 10515 1505 10555
rect 1435 10475 1505 10515
rect 1435 10435 1450 10475
rect 1490 10435 1505 10475
rect 1435 10395 1505 10435
rect 1435 10355 1450 10395
rect 1490 10355 1505 10395
rect 1435 10315 1505 10355
rect 1435 10275 1450 10315
rect 1490 10275 1505 10315
rect 1435 10260 1505 10275
rect 1550 12235 1620 12255
rect 1550 12195 1565 12235
rect 1605 12195 1620 12235
rect 1550 12155 1620 12195
rect 1550 12115 1565 12155
rect 1605 12115 1620 12155
rect 1550 12075 1620 12115
rect 1550 12035 1565 12075
rect 1605 12035 1620 12075
rect 1550 11995 1620 12035
rect 1550 11955 1565 11995
rect 1605 11955 1620 11995
rect 1550 11915 1620 11955
rect 1550 11875 1565 11915
rect 1605 11875 1620 11915
rect 1550 11835 1620 11875
rect 1550 11795 1565 11835
rect 1605 11795 1620 11835
rect 1550 11755 1620 11795
rect 1550 11715 1565 11755
rect 1605 11715 1620 11755
rect 1550 11675 1620 11715
rect 1550 11635 1565 11675
rect 1605 11635 1620 11675
rect 1550 11595 1620 11635
rect 1550 11555 1565 11595
rect 1605 11555 1620 11595
rect 1550 11515 1620 11555
rect 1550 11475 1565 11515
rect 1605 11475 1620 11515
rect 1550 11435 1620 11475
rect 1550 11395 1565 11435
rect 1605 11395 1620 11435
rect 1550 11355 1620 11395
rect 1550 11315 1565 11355
rect 1605 11315 1620 11355
rect 1550 11275 1620 11315
rect 1550 11235 1565 11275
rect 1605 11235 1620 11275
rect 1550 11195 1620 11235
rect 1550 11155 1565 11195
rect 1605 11155 1620 11195
rect 1550 11115 1620 11155
rect 1550 11075 1565 11115
rect 1605 11075 1620 11115
rect 1550 11035 1620 11075
rect 1550 10995 1565 11035
rect 1605 10995 1620 11035
rect 1550 10955 1620 10995
rect 1550 10915 1565 10955
rect 1605 10915 1620 10955
rect 1550 10875 1620 10915
rect 1550 10835 1565 10875
rect 1605 10835 1620 10875
rect 1550 10795 1620 10835
rect 1550 10755 1565 10795
rect 1605 10755 1620 10795
rect 1550 10715 1620 10755
rect 1550 10675 1565 10715
rect 1605 10675 1620 10715
rect 1550 10635 1620 10675
rect 1550 10595 1565 10635
rect 1605 10595 1620 10635
rect 1550 10555 1620 10595
rect 1550 10515 1565 10555
rect 1605 10515 1620 10555
rect 1550 10475 1620 10515
rect 1550 10435 1565 10475
rect 1605 10435 1620 10475
rect 1550 10395 1620 10435
rect 1550 10355 1565 10395
rect 1605 10355 1620 10395
rect 1550 10315 1620 10355
rect 1550 10275 1565 10315
rect 1605 10275 1620 10315
rect 1550 10150 1620 10275
rect 1665 12235 1735 12340
rect 1665 12195 1680 12235
rect 1720 12195 1735 12235
rect 1665 12155 1735 12195
rect 1665 12115 1680 12155
rect 1720 12115 1735 12155
rect 1665 12075 1735 12115
rect 1665 12035 1680 12075
rect 1720 12035 1735 12075
rect 1665 11995 1735 12035
rect 1665 11955 1680 11995
rect 1720 11955 1735 11995
rect 1665 11915 1735 11955
rect 1665 11875 1680 11915
rect 1720 11875 1735 11915
rect 1665 11835 1735 11875
rect 1665 11795 1680 11835
rect 1720 11795 1735 11835
rect 1665 11755 1735 11795
rect 1665 11715 1680 11755
rect 1720 11715 1735 11755
rect 1665 11675 1735 11715
rect 1665 11635 1680 11675
rect 1720 11635 1735 11675
rect 1665 11595 1735 11635
rect 1665 11555 1680 11595
rect 1720 11555 1735 11595
rect 1665 11515 1735 11555
rect 1665 11475 1680 11515
rect 1720 11475 1735 11515
rect 1665 11435 1735 11475
rect 1665 11395 1680 11435
rect 1720 11395 1735 11435
rect 1665 11355 1735 11395
rect 1665 11315 1680 11355
rect 1720 11315 1735 11355
rect 1665 11275 1735 11315
rect 1665 11235 1680 11275
rect 1720 11235 1735 11275
rect 1665 11195 1735 11235
rect 1665 11155 1680 11195
rect 1720 11155 1735 11195
rect 1665 11115 1735 11155
rect 1665 11075 1680 11115
rect 1720 11075 1735 11115
rect 1665 11035 1735 11075
rect 1665 10995 1680 11035
rect 1720 10995 1735 11035
rect 1665 10955 1735 10995
rect 1665 10915 1680 10955
rect 1720 10915 1735 10955
rect 1665 10875 1735 10915
rect 1665 10835 1680 10875
rect 1720 10835 1735 10875
rect 1665 10795 1735 10835
rect 1665 10755 1680 10795
rect 1720 10755 1735 10795
rect 1665 10715 1735 10755
rect 1665 10675 1680 10715
rect 1720 10675 1735 10715
rect 1665 10635 1735 10675
rect 1665 10595 1680 10635
rect 1720 10595 1735 10635
rect 1665 10555 1735 10595
rect 1665 10515 1680 10555
rect 1720 10515 1735 10555
rect 1665 10475 1735 10515
rect 1665 10435 1680 10475
rect 1720 10435 1735 10475
rect 1665 10395 1735 10435
rect 1665 10355 1680 10395
rect 1720 10355 1735 10395
rect 1665 10315 1735 10355
rect 1665 10275 1680 10315
rect 1720 10275 1735 10315
rect 1665 10260 1735 10275
rect 1780 12235 1850 12255
rect 1780 12195 1795 12235
rect 1835 12195 1850 12235
rect 1780 12155 1850 12195
rect 1780 12115 1795 12155
rect 1835 12115 1850 12155
rect 1780 12075 1850 12115
rect 1780 12035 1795 12075
rect 1835 12035 1850 12075
rect 1780 11995 1850 12035
rect 1780 11955 1795 11995
rect 1835 11955 1850 11995
rect 1780 11915 1850 11955
rect 1780 11875 1795 11915
rect 1835 11875 1850 11915
rect 1780 11835 1850 11875
rect 1780 11795 1795 11835
rect 1835 11795 1850 11835
rect 1780 11755 1850 11795
rect 1780 11715 1795 11755
rect 1835 11715 1850 11755
rect 1780 11675 1850 11715
rect 1780 11635 1795 11675
rect 1835 11635 1850 11675
rect 1780 11595 1850 11635
rect 1780 11555 1795 11595
rect 1835 11555 1850 11595
rect 1780 11515 1850 11555
rect 1780 11475 1795 11515
rect 1835 11475 1850 11515
rect 1780 11435 1850 11475
rect 1780 11395 1795 11435
rect 1835 11395 1850 11435
rect 1780 11355 1850 11395
rect 1780 11315 1795 11355
rect 1835 11315 1850 11355
rect 1780 11275 1850 11315
rect 1780 11235 1795 11275
rect 1835 11235 1850 11275
rect 1780 11195 1850 11235
rect 1780 11155 1795 11195
rect 1835 11155 1850 11195
rect 1780 11115 1850 11155
rect 1780 11075 1795 11115
rect 1835 11075 1850 11115
rect 1780 11035 1850 11075
rect 1780 10995 1795 11035
rect 1835 10995 1850 11035
rect 1780 10955 1850 10995
rect 1780 10915 1795 10955
rect 1835 10915 1850 10955
rect 1780 10875 1850 10915
rect 1780 10835 1795 10875
rect 1835 10835 1850 10875
rect 1780 10795 1850 10835
rect 1780 10755 1795 10795
rect 1835 10755 1850 10795
rect 1780 10715 1850 10755
rect 1780 10675 1795 10715
rect 1835 10675 1850 10715
rect 1780 10635 1850 10675
rect 1780 10595 1795 10635
rect 1835 10595 1850 10635
rect 1780 10555 1850 10595
rect 1780 10515 1795 10555
rect 1835 10515 1850 10555
rect 1780 10475 1850 10515
rect 1780 10435 1795 10475
rect 1835 10435 1850 10475
rect 1780 10395 1850 10435
rect 1780 10355 1795 10395
rect 1835 10355 1850 10395
rect 1780 10315 1850 10355
rect 1780 10275 1795 10315
rect 1835 10275 1850 10315
rect 1780 10150 1850 10275
rect 1895 12235 1965 12340
rect 1895 12195 1910 12235
rect 1950 12195 1965 12235
rect 1895 12155 1965 12195
rect 1895 12115 1910 12155
rect 1950 12115 1965 12155
rect 1895 12075 1965 12115
rect 1895 12035 1910 12075
rect 1950 12035 1965 12075
rect 1895 11995 1965 12035
rect 1895 11955 1910 11995
rect 1950 11955 1965 11995
rect 1895 11915 1965 11955
rect 1895 11875 1910 11915
rect 1950 11875 1965 11915
rect 1895 11835 1965 11875
rect 1895 11795 1910 11835
rect 1950 11795 1965 11835
rect 1895 11755 1965 11795
rect 1895 11715 1910 11755
rect 1950 11715 1965 11755
rect 1895 11675 1965 11715
rect 1895 11635 1910 11675
rect 1950 11635 1965 11675
rect 1895 11595 1965 11635
rect 1895 11555 1910 11595
rect 1950 11555 1965 11595
rect 1895 11515 1965 11555
rect 1895 11475 1910 11515
rect 1950 11475 1965 11515
rect 1895 11435 1965 11475
rect 1895 11395 1910 11435
rect 1950 11395 1965 11435
rect 1895 11355 1965 11395
rect 1895 11315 1910 11355
rect 1950 11315 1965 11355
rect 1895 11275 1965 11315
rect 1895 11235 1910 11275
rect 1950 11235 1965 11275
rect 1895 11195 1965 11235
rect 1895 11155 1910 11195
rect 1950 11155 1965 11195
rect 1895 11115 1965 11155
rect 1895 11075 1910 11115
rect 1950 11075 1965 11115
rect 1895 11035 1965 11075
rect 1895 10995 1910 11035
rect 1950 10995 1965 11035
rect 1895 10955 1965 10995
rect 1895 10915 1910 10955
rect 1950 10915 1965 10955
rect 1895 10875 1965 10915
rect 1895 10835 1910 10875
rect 1950 10835 1965 10875
rect 1895 10795 1965 10835
rect 1895 10755 1910 10795
rect 1950 10755 1965 10795
rect 1895 10715 1965 10755
rect 1895 10675 1910 10715
rect 1950 10675 1965 10715
rect 1895 10635 1965 10675
rect 1895 10595 1910 10635
rect 1950 10595 1965 10635
rect 1895 10555 1965 10595
rect 1895 10515 1910 10555
rect 1950 10515 1965 10555
rect 1895 10475 1965 10515
rect 1895 10435 1910 10475
rect 1950 10435 1965 10475
rect 1895 10395 1965 10435
rect 1895 10355 1910 10395
rect 1950 10355 1965 10395
rect 1895 10315 1965 10355
rect 1895 10275 1910 10315
rect 1950 10275 1965 10315
rect 1895 10260 1965 10275
rect 2010 12235 2080 12255
rect 2010 12195 2025 12235
rect 2065 12195 2080 12235
rect 2010 12155 2080 12195
rect 2010 12115 2025 12155
rect 2065 12115 2080 12155
rect 2010 12075 2080 12115
rect 2010 12035 2025 12075
rect 2065 12035 2080 12075
rect 2010 11995 2080 12035
rect 2010 11955 2025 11995
rect 2065 11955 2080 11995
rect 2010 11915 2080 11955
rect 2010 11875 2025 11915
rect 2065 11875 2080 11915
rect 2010 11835 2080 11875
rect 2010 11795 2025 11835
rect 2065 11795 2080 11835
rect 2010 11755 2080 11795
rect 2010 11715 2025 11755
rect 2065 11715 2080 11755
rect 2010 11675 2080 11715
rect 2010 11635 2025 11675
rect 2065 11635 2080 11675
rect 2010 11595 2080 11635
rect 2010 11555 2025 11595
rect 2065 11555 2080 11595
rect 2010 11515 2080 11555
rect 2010 11475 2025 11515
rect 2065 11475 2080 11515
rect 2010 11435 2080 11475
rect 2010 11395 2025 11435
rect 2065 11395 2080 11435
rect 2010 11355 2080 11395
rect 2010 11315 2025 11355
rect 2065 11315 2080 11355
rect 2010 11275 2080 11315
rect 2010 11235 2025 11275
rect 2065 11235 2080 11275
rect 2010 11195 2080 11235
rect 2010 11155 2025 11195
rect 2065 11155 2080 11195
rect 2010 11115 2080 11155
rect 2010 11075 2025 11115
rect 2065 11075 2080 11115
rect 2010 11035 2080 11075
rect 2010 10995 2025 11035
rect 2065 10995 2080 11035
rect 2010 10955 2080 10995
rect 2010 10915 2025 10955
rect 2065 10915 2080 10955
rect 2010 10875 2080 10915
rect 2010 10835 2025 10875
rect 2065 10835 2080 10875
rect 2010 10795 2080 10835
rect 2010 10755 2025 10795
rect 2065 10755 2080 10795
rect 2010 10715 2080 10755
rect 2010 10675 2025 10715
rect 2065 10675 2080 10715
rect 2010 10635 2080 10675
rect 2010 10595 2025 10635
rect 2065 10595 2080 10635
rect 2010 10555 2080 10595
rect 2010 10515 2025 10555
rect 2065 10515 2080 10555
rect 2010 10475 2080 10515
rect 2010 10435 2025 10475
rect 2065 10435 2080 10475
rect 2010 10395 2080 10435
rect 2010 10355 2025 10395
rect 2065 10355 2080 10395
rect 2010 10315 2080 10355
rect 2010 10275 2025 10315
rect 2065 10275 2080 10315
rect 2010 10150 2080 10275
rect 2125 12235 2195 12340
rect 2125 12195 2140 12235
rect 2180 12195 2195 12235
rect 2125 12155 2195 12195
rect 2125 12115 2140 12155
rect 2180 12115 2195 12155
rect 2125 12075 2195 12115
rect 2125 12035 2140 12075
rect 2180 12035 2195 12075
rect 2125 11995 2195 12035
rect 2125 11955 2140 11995
rect 2180 11955 2195 11995
rect 2125 11915 2195 11955
rect 2125 11875 2140 11915
rect 2180 11875 2195 11915
rect 2125 11835 2195 11875
rect 2125 11795 2140 11835
rect 2180 11795 2195 11835
rect 2125 11755 2195 11795
rect 2125 11715 2140 11755
rect 2180 11715 2195 11755
rect 2125 11675 2195 11715
rect 2125 11635 2140 11675
rect 2180 11635 2195 11675
rect 2125 11595 2195 11635
rect 2125 11555 2140 11595
rect 2180 11555 2195 11595
rect 2125 11515 2195 11555
rect 2125 11475 2140 11515
rect 2180 11475 2195 11515
rect 2125 11435 2195 11475
rect 2125 11395 2140 11435
rect 2180 11395 2195 11435
rect 2125 11355 2195 11395
rect 2125 11315 2140 11355
rect 2180 11315 2195 11355
rect 2125 11275 2195 11315
rect 2125 11235 2140 11275
rect 2180 11235 2195 11275
rect 2125 11195 2195 11235
rect 2125 11155 2140 11195
rect 2180 11155 2195 11195
rect 2125 11115 2195 11155
rect 2125 11075 2140 11115
rect 2180 11075 2195 11115
rect 2125 11035 2195 11075
rect 2125 10995 2140 11035
rect 2180 10995 2195 11035
rect 2125 10955 2195 10995
rect 2125 10915 2140 10955
rect 2180 10915 2195 10955
rect 2125 10875 2195 10915
rect 2125 10835 2140 10875
rect 2180 10835 2195 10875
rect 2125 10795 2195 10835
rect 2125 10755 2140 10795
rect 2180 10755 2195 10795
rect 2125 10715 2195 10755
rect 2125 10675 2140 10715
rect 2180 10675 2195 10715
rect 2125 10635 2195 10675
rect 2125 10595 2140 10635
rect 2180 10595 2195 10635
rect 2125 10555 2195 10595
rect 2125 10515 2140 10555
rect 2180 10515 2195 10555
rect 2125 10475 2195 10515
rect 2125 10435 2140 10475
rect 2180 10435 2195 10475
rect 2125 10395 2195 10435
rect 2125 10355 2140 10395
rect 2180 10355 2195 10395
rect 2125 10315 2195 10355
rect 2125 10275 2140 10315
rect 2180 10275 2195 10315
rect 2125 10260 2195 10275
rect 2240 12235 2310 12255
rect 2240 12195 2255 12235
rect 2295 12195 2310 12235
rect 2240 12155 2310 12195
rect 2240 12115 2255 12155
rect 2295 12115 2310 12155
rect 2240 12075 2310 12115
rect 2240 12035 2255 12075
rect 2295 12035 2310 12075
rect 2240 11995 2310 12035
rect 2240 11955 2255 11995
rect 2295 11955 2310 11995
rect 2240 11915 2310 11955
rect 2240 11875 2255 11915
rect 2295 11875 2310 11915
rect 2240 11835 2310 11875
rect 2240 11795 2255 11835
rect 2295 11795 2310 11835
rect 2240 11755 2310 11795
rect 2240 11715 2255 11755
rect 2295 11715 2310 11755
rect 2240 11675 2310 11715
rect 2240 11635 2255 11675
rect 2295 11635 2310 11675
rect 2240 11595 2310 11635
rect 2240 11555 2255 11595
rect 2295 11555 2310 11595
rect 2240 11515 2310 11555
rect 2240 11475 2255 11515
rect 2295 11475 2310 11515
rect 2240 11435 2310 11475
rect 2240 11395 2255 11435
rect 2295 11395 2310 11435
rect 2240 11355 2310 11395
rect 2240 11315 2255 11355
rect 2295 11315 2310 11355
rect 2240 11275 2310 11315
rect 2240 11235 2255 11275
rect 2295 11235 2310 11275
rect 2240 11195 2310 11235
rect 2240 11155 2255 11195
rect 2295 11155 2310 11195
rect 2240 11115 2310 11155
rect 2240 11075 2255 11115
rect 2295 11075 2310 11115
rect 2240 11035 2310 11075
rect 2240 10995 2255 11035
rect 2295 10995 2310 11035
rect 2240 10955 2310 10995
rect 2240 10915 2255 10955
rect 2295 10915 2310 10955
rect 2240 10875 2310 10915
rect 2240 10835 2255 10875
rect 2295 10835 2310 10875
rect 2240 10795 2310 10835
rect 2240 10755 2255 10795
rect 2295 10755 2310 10795
rect 2240 10715 2310 10755
rect 2240 10675 2255 10715
rect 2295 10675 2310 10715
rect 2240 10635 2310 10675
rect 2240 10595 2255 10635
rect 2295 10595 2310 10635
rect 2240 10555 2310 10595
rect 2240 10515 2255 10555
rect 2295 10515 2310 10555
rect 2240 10475 2310 10515
rect 2240 10435 2255 10475
rect 2295 10435 2310 10475
rect 2240 10395 2310 10435
rect 2240 10355 2255 10395
rect 2295 10355 2310 10395
rect 2240 10315 2310 10355
rect 2240 10275 2255 10315
rect 2295 10275 2310 10315
rect 2240 10150 2310 10275
rect 2355 12235 2425 12340
rect 2355 12195 2370 12235
rect 2410 12195 2425 12235
rect 2355 12155 2425 12195
rect 2355 12115 2370 12155
rect 2410 12115 2425 12155
rect 2355 12075 2425 12115
rect 2355 12035 2370 12075
rect 2410 12035 2425 12075
rect 2355 11995 2425 12035
rect 2355 11955 2370 11995
rect 2410 11955 2425 11995
rect 2355 11915 2425 11955
rect 2355 11875 2370 11915
rect 2410 11875 2425 11915
rect 2355 11835 2425 11875
rect 2355 11795 2370 11835
rect 2410 11795 2425 11835
rect 2355 11755 2425 11795
rect 2355 11715 2370 11755
rect 2410 11715 2425 11755
rect 2355 11675 2425 11715
rect 2355 11635 2370 11675
rect 2410 11635 2425 11675
rect 2355 11595 2425 11635
rect 2355 11555 2370 11595
rect 2410 11555 2425 11595
rect 2355 11515 2425 11555
rect 2355 11475 2370 11515
rect 2410 11475 2425 11515
rect 2355 11435 2425 11475
rect 2355 11395 2370 11435
rect 2410 11395 2425 11435
rect 2355 11355 2425 11395
rect 2355 11315 2370 11355
rect 2410 11315 2425 11355
rect 2355 11275 2425 11315
rect 2355 11235 2370 11275
rect 2410 11235 2425 11275
rect 2355 11195 2425 11235
rect 2355 11155 2370 11195
rect 2410 11155 2425 11195
rect 2355 11115 2425 11155
rect 2355 11075 2370 11115
rect 2410 11075 2425 11115
rect 2355 11035 2425 11075
rect 2355 10995 2370 11035
rect 2410 10995 2425 11035
rect 2355 10955 2425 10995
rect 2355 10915 2370 10955
rect 2410 10915 2425 10955
rect 2355 10875 2425 10915
rect 2355 10835 2370 10875
rect 2410 10835 2425 10875
rect 2355 10795 2425 10835
rect 2355 10755 2370 10795
rect 2410 10755 2425 10795
rect 2355 10715 2425 10755
rect 2355 10675 2370 10715
rect 2410 10675 2425 10715
rect 2355 10635 2425 10675
rect 2355 10595 2370 10635
rect 2410 10595 2425 10635
rect 2355 10555 2425 10595
rect 2355 10515 2370 10555
rect 2410 10515 2425 10555
rect 2355 10475 2425 10515
rect 2355 10435 2370 10475
rect 2410 10435 2425 10475
rect 2355 10395 2425 10435
rect 2355 10355 2370 10395
rect 2410 10355 2425 10395
rect 2355 10315 2425 10355
rect 2355 10275 2370 10315
rect 2410 10275 2425 10315
rect 2355 10260 2425 10275
rect 2470 12235 2540 12255
rect 2470 12195 2485 12235
rect 2525 12195 2540 12235
rect 2470 12155 2540 12195
rect 2470 12115 2485 12155
rect 2525 12115 2540 12155
rect 2470 12075 2540 12115
rect 2470 12035 2485 12075
rect 2525 12035 2540 12075
rect 2470 11995 2540 12035
rect 2470 11955 2485 11995
rect 2525 11955 2540 11995
rect 2470 11915 2540 11955
rect 2470 11875 2485 11915
rect 2525 11875 2540 11915
rect 2470 11835 2540 11875
rect 2470 11795 2485 11835
rect 2525 11795 2540 11835
rect 2470 11755 2540 11795
rect 2470 11715 2485 11755
rect 2525 11715 2540 11755
rect 2470 11675 2540 11715
rect 2470 11635 2485 11675
rect 2525 11635 2540 11675
rect 2470 11595 2540 11635
rect 2470 11555 2485 11595
rect 2525 11555 2540 11595
rect 2470 11515 2540 11555
rect 2470 11475 2485 11515
rect 2525 11475 2540 11515
rect 2470 11435 2540 11475
rect 2470 11395 2485 11435
rect 2525 11395 2540 11435
rect 2470 11355 2540 11395
rect 2470 11315 2485 11355
rect 2525 11315 2540 11355
rect 2470 11275 2540 11315
rect 2470 11235 2485 11275
rect 2525 11235 2540 11275
rect 2470 11195 2540 11235
rect 2470 11155 2485 11195
rect 2525 11155 2540 11195
rect 2470 11115 2540 11155
rect 2470 11075 2485 11115
rect 2525 11075 2540 11115
rect 2470 11035 2540 11075
rect 2470 10995 2485 11035
rect 2525 10995 2540 11035
rect 2470 10955 2540 10995
rect 2470 10915 2485 10955
rect 2525 10915 2540 10955
rect 2470 10875 2540 10915
rect 2470 10835 2485 10875
rect 2525 10835 2540 10875
rect 2470 10795 2540 10835
rect 2470 10755 2485 10795
rect 2525 10755 2540 10795
rect 2470 10715 2540 10755
rect 2470 10675 2485 10715
rect 2525 10675 2540 10715
rect 2470 10635 2540 10675
rect 2470 10595 2485 10635
rect 2525 10595 2540 10635
rect 2470 10555 2540 10595
rect 2470 10515 2485 10555
rect 2525 10515 2540 10555
rect 2470 10475 2540 10515
rect 2470 10435 2485 10475
rect 2525 10435 2540 10475
rect 2470 10395 2540 10435
rect 2470 10355 2485 10395
rect 2525 10355 2540 10395
rect 2470 10315 2540 10355
rect 2470 10275 2485 10315
rect 2525 10275 2540 10315
rect 2470 10150 2540 10275
rect 2655 12155 2755 12285
rect 2655 12115 2685 12155
rect 2725 12115 2755 12155
rect 2655 11995 2755 12115
rect 2655 11955 2685 11995
rect 2725 11955 2755 11995
rect 2655 11835 2755 11955
rect 2655 11795 2685 11835
rect 2725 11795 2755 11835
rect 2655 11675 2755 11795
rect 2655 11635 2685 11675
rect 2725 11635 2755 11675
rect 2655 11515 2755 11635
rect 2655 11475 2685 11515
rect 2725 11475 2755 11515
rect 2655 11355 2755 11475
rect 2655 11315 2685 11355
rect 2725 11315 2755 11355
rect 2655 11195 2755 11315
rect 2655 11155 2685 11195
rect 2725 11155 2755 11195
rect 2655 10955 2755 11155
rect 2655 10915 2685 10955
rect 2725 10915 2755 10955
rect 2655 10795 2755 10915
rect 2655 10755 2685 10795
rect 2725 10755 2755 10795
rect 2655 10635 2755 10755
rect 2655 10595 2685 10635
rect 2725 10595 2755 10635
rect 2655 10475 2755 10595
rect 2655 10435 2685 10475
rect 2725 10435 2755 10475
rect 2655 10315 2755 10435
rect 2655 10275 2685 10315
rect 2725 10275 2755 10315
rect 2655 10230 2755 10275
rect -1050 10120 3300 10150
rect -620 10030 880 10060
rect -620 9990 -390 10030
rect -350 9990 -230 10030
rect -190 9990 -70 10030
rect -30 9990 90 10030
rect 130 9990 250 10030
rect 290 9990 410 10030
rect 450 9990 570 10030
rect 610 9990 730 10030
rect 770 9990 880 10030
rect -620 9960 880 9990
rect 1260 10030 2755 10060
rect 1260 9990 1290 10030
rect 1330 9990 1450 10030
rect 1490 9990 1610 10030
rect 1650 9990 1770 10030
rect 1810 9990 1930 10030
rect 1970 9990 2090 10030
rect 2130 9990 2250 10030
rect 2290 9990 2410 10030
rect 2450 9990 2755 10030
rect 1260 9960 2755 9990
<< end >>
