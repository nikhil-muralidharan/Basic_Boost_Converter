magic
tech sky130A
timestamp 1638706231
<< end >>
