magic
tech sky130A
timestamp 1659419658
<< nwell >>
rect -180 170 485 330
<< pmoslvt >>
rect 0 200 35 300
rect 85 200 120 300
rect 330 200 365 300
<< nmoslvt >>
rect 0 5 15 105
rect 65 5 80 105
rect 330 5 345 105
<< ndiff >>
rect -50 90 0 105
rect -50 20 -35 90
rect -15 20 0 90
rect -50 5 0 20
rect 15 90 65 105
rect 15 20 30 90
rect 50 20 65 90
rect 15 5 65 20
rect 80 90 130 105
rect 80 20 95 90
rect 115 20 130 90
rect 80 5 130 20
rect 280 90 330 105
rect 280 20 295 90
rect 315 20 330 90
rect 280 5 330 20
rect 345 90 395 105
rect 345 20 360 90
rect 380 20 395 90
rect 345 5 395 20
<< pdiff >>
rect -50 285 0 300
rect -50 215 -35 285
rect -15 215 0 285
rect -50 200 0 215
rect 35 285 85 300
rect 35 215 50 285
rect 70 215 85 285
rect 35 200 85 215
rect 120 285 170 300
rect 120 215 135 285
rect 155 215 170 285
rect 120 200 170 215
rect 280 285 330 300
rect 280 215 295 285
rect 315 215 330 285
rect 280 200 330 215
rect 365 285 415 300
rect 365 215 380 285
rect 400 215 415 285
rect 365 200 415 215
<< ndiffc >>
rect -35 20 -15 90
rect 30 20 50 90
rect 95 20 115 90
rect 295 20 315 90
rect 360 20 380 90
<< pdiffc >>
rect -35 215 -15 285
rect 50 215 70 285
rect 135 215 155 285
rect 295 215 315 285
rect 380 215 400 285
<< psubdiff >>
rect -130 90 -80 105
rect -130 20 -115 90
rect -95 20 -80 90
rect -130 5 -80 20
<< nsubdiff >>
rect -130 285 -80 300
rect -130 215 -115 285
rect -95 215 -80 285
rect -130 200 -80 215
<< psubdiffcont >>
rect -115 20 -95 90
<< nsubdiffcont >>
rect -115 215 -95 285
<< poly >>
rect -5 380 35 390
rect -5 360 5 380
rect 25 360 35 380
rect -5 350 35 360
rect 0 300 35 350
rect 85 380 125 390
rect 85 360 95 380
rect 115 360 125 380
rect 85 350 125 360
rect 330 370 370 380
rect 330 350 340 370
rect 360 350 370 370
rect 85 300 120 350
rect 330 340 370 350
rect 330 300 365 340
rect 0 185 35 200
rect 85 185 120 200
rect 330 185 365 200
rect 0 105 15 120
rect 65 105 80 120
rect 330 105 345 185
rect 0 -80 15 5
rect -25 -90 15 -80
rect -25 -110 -15 -90
rect 5 -110 15 -90
rect -25 -120 15 -110
rect 65 -80 80 5
rect 330 -30 345 5
rect 330 -40 370 -30
rect 330 -60 340 -40
rect 360 -60 370 -40
rect 330 -70 370 -60
rect 65 -90 105 -80
rect 65 -110 75 -90
rect 95 -110 105 -90
rect 65 -120 105 -110
<< polycont >>
rect 5 360 25 380
rect 95 360 115 380
rect 340 350 360 370
rect -15 -110 5 -90
rect 340 -60 360 -40
rect 75 -110 95 -90
<< locali >>
rect -180 410 360 430
rect 10 390 30 410
rect -5 380 35 390
rect -5 360 5 380
rect 25 360 35 380
rect -5 350 35 360
rect 85 380 125 390
rect 340 380 360 410
rect 85 360 95 380
rect 115 375 125 380
rect 115 360 240 375
rect 85 350 240 360
rect -125 285 -85 295
rect -125 215 -115 285
rect -95 215 -85 285
rect -125 205 -85 215
rect -45 285 -5 295
rect -45 215 -35 285
rect -15 215 -5 285
rect -45 205 -5 215
rect 40 285 80 295
rect 40 215 50 285
rect 70 215 80 285
rect 40 205 80 215
rect 125 285 165 295
rect 125 215 135 285
rect 155 215 165 285
rect 125 205 165 215
rect -35 100 -15 205
rect 50 180 70 205
rect 30 170 75 180
rect 30 140 40 170
rect 70 140 75 170
rect 135 140 155 205
rect 30 130 75 140
rect 30 100 50 130
rect 95 120 155 140
rect 220 160 240 350
rect 330 370 370 380
rect 330 350 340 370
rect 360 350 370 370
rect 330 340 370 350
rect 285 285 325 295
rect 285 215 295 285
rect 315 215 325 285
rect 285 205 325 215
rect 370 285 410 295
rect 370 215 380 285
rect 400 215 410 285
rect 370 205 410 215
rect 295 160 315 205
rect 220 140 315 160
rect 95 100 115 120
rect -125 90 -85 100
rect -125 20 -115 90
rect -95 20 -85 90
rect -125 10 -85 20
rect -45 90 -5 100
rect -45 20 -35 90
rect -15 20 -5 90
rect -45 -15 -5 20
rect 20 90 60 100
rect 20 20 30 90
rect 50 20 60 90
rect 20 10 60 20
rect 85 90 125 100
rect 85 20 95 90
rect 115 20 125 90
rect -45 -35 -35 -15
rect -15 -35 -5 -15
rect -45 -45 -5 -35
rect 85 -15 125 20
rect 85 -35 95 -15
rect 115 -35 125 -15
rect 85 -45 125 -35
rect -25 -90 15 -80
rect -25 -110 -15 -90
rect 5 -110 15 -90
rect -25 -120 15 -110
rect 65 -90 105 -80
rect 220 -90 240 140
rect 295 100 315 140
rect 285 90 325 100
rect 285 20 295 90
rect 315 20 325 90
rect 285 10 325 20
rect 350 90 390 100
rect 350 20 360 90
rect 380 20 390 90
rect 350 10 390 20
rect 330 -40 370 -30
rect 330 -60 340 -40
rect 360 -60 370 -40
rect 330 -70 370 -60
rect 65 -110 75 -90
rect 95 -110 240 -90
rect 65 -120 105 -110
rect -5 -140 15 -120
rect 340 -140 360 -70
rect -5 -160 360 -140
<< viali >>
rect -115 215 -95 285
rect 40 140 70 170
rect 380 215 400 285
rect -115 20 -95 90
rect -35 -35 -15 -15
rect 95 -35 115 -15
rect 360 20 380 90
<< metal1 >>
rect -180 285 485 295
rect -180 215 -115 285
rect -95 215 380 285
rect 400 215 485 285
rect -180 205 485 215
rect 30 170 75 180
rect 30 140 40 170
rect 70 140 75 170
rect 30 130 75 140
rect -175 90 485 100
rect -175 20 -115 90
rect -95 20 360 90
rect 380 20 485 90
rect -175 10 485 20
rect -45 -15 -5 -5
rect -45 -35 -35 -15
rect -15 -35 -5 -15
rect -45 -190 -5 -35
rect 85 -15 125 -5
rect 85 -35 95 -15
rect 115 -35 125 -15
rect 85 -190 125 -35
<< via1 >>
rect 40 140 70 170
<< metal2 >>
rect 45 180 75 500
rect 30 170 75 180
rect 30 140 40 170
rect 70 140 75 170
rect 30 130 75 140
<< labels >>
rlabel metal1 -180 250 -180 250 7 VP
port 1 w
rlabel metal1 -175 50 -175 50 7 VN
port 2 w
rlabel metal1 -25 -190 -25 -190 5 IN1
port 3 s
rlabel metal1 105 -190 105 -190 5 IN2
port 4 s
rlabel locali -180 420 -180 420 7 S
port 5 w
rlabel metal2 60 500 60 500 1 Y
port 6 n
<< end >>
