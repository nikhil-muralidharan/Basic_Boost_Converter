magic
tech sky130A
timestamp 1640179548
<< error_p >>
rect -333 12270 -320 12283
rect -345 10245 -320 12270
rect -333 10232 -320 10245
<< nmos >>
rect -320 10245 -305 12270
<< ndiff >>
rect -305 12235 -205 12270
rect -305 12195 -275 12235
rect -235 12195 -205 12235
rect -305 12155 -205 12195
rect -305 12115 -275 12155
rect -235 12115 -205 12155
rect -305 12075 -205 12115
rect -305 12035 -275 12075
rect -235 12035 -205 12075
rect -305 11995 -205 12035
rect -305 11955 -275 11995
rect -235 11955 -205 11995
rect -305 11915 -205 11955
rect -305 11875 -275 11915
rect -235 11875 -205 11915
rect -305 11835 -205 11875
rect -305 11795 -275 11835
rect -235 11795 -205 11835
rect -305 11755 -205 11795
rect -305 11715 -275 11755
rect -235 11715 -205 11755
rect -305 11675 -205 11715
rect -305 11635 -275 11675
rect -235 11635 -205 11675
rect -305 11595 -205 11635
rect -305 11555 -275 11595
rect -235 11555 -205 11595
rect -305 11515 -205 11555
rect -305 11475 -275 11515
rect -235 11475 -205 11515
rect -305 11435 -205 11475
rect -305 11395 -275 11435
rect -235 11395 -205 11435
rect -305 11355 -205 11395
rect -305 11315 -275 11355
rect -235 11315 -205 11355
rect -305 11275 -205 11315
rect -305 11235 -275 11275
rect -235 11235 -205 11275
rect -305 11195 -205 11235
rect -305 11155 -275 11195
rect -235 11155 -205 11195
rect -305 11115 -205 11155
rect -305 11075 -275 11115
rect -235 11075 -205 11115
rect -305 11035 -205 11075
rect -305 10995 -275 11035
rect -235 10995 -205 11035
rect -305 10955 -205 10995
rect -305 10915 -275 10955
rect -235 10915 -205 10955
rect -305 10875 -205 10915
rect -305 10835 -275 10875
rect -235 10835 -205 10875
rect -305 10795 -205 10835
rect -305 10755 -275 10795
rect -235 10755 -205 10795
rect -305 10715 -205 10755
rect -305 10675 -275 10715
rect -235 10675 -205 10715
rect -305 10635 -205 10675
rect -305 10595 -275 10635
rect -235 10595 -205 10635
rect -305 10555 -205 10595
rect -305 10515 -275 10555
rect -235 10515 -205 10555
rect -305 10475 -205 10515
rect -305 10435 -275 10475
rect -235 10435 -205 10475
rect -305 10395 -205 10435
rect -305 10355 -275 10395
rect -235 10355 -205 10395
rect -305 10315 -205 10355
rect -305 10275 -275 10315
rect -235 10275 -205 10315
rect -305 10245 -205 10275
<< ndiffc >>
rect -275 12195 -235 12235
rect -275 12115 -235 12155
rect -275 12035 -235 12075
rect -275 11955 -235 11995
rect -275 11875 -235 11915
rect -275 11795 -235 11835
rect -275 11715 -235 11755
rect -275 11635 -235 11675
rect -275 11555 -235 11595
rect -275 11475 -235 11515
rect -275 11395 -235 11435
rect -275 11315 -235 11355
rect -275 11235 -235 11275
rect -275 11155 -235 11195
rect -275 11075 -235 11115
rect -275 10995 -235 11035
rect -275 10915 -235 10955
rect -275 10835 -235 10875
rect -275 10755 -235 10795
rect -275 10675 -235 10715
rect -275 10595 -235 10635
rect -275 10515 -235 10555
rect -275 10435 -235 10475
rect -275 10355 -235 10395
rect -275 10275 -235 10315
<< poly >>
rect -320 12270 -305 12290
rect -320 10170 -305 10245
rect -345 10160 -305 10170
rect -345 10140 -335 10160
rect -315 10140 -305 10160
rect -345 10130 -305 10140
<< polycont >>
rect -335 10140 -315 10160
<< locali >>
rect -290 12235 -220 12255
rect -290 12195 -275 12235
rect -235 12195 -220 12235
rect -290 12155 -220 12195
rect -290 12115 -275 12155
rect -235 12115 -220 12155
rect -290 12075 -220 12115
rect -290 12035 -275 12075
rect -235 12035 -220 12075
rect -290 11995 -220 12035
rect -290 11955 -275 11995
rect -235 11955 -220 11995
rect -290 11915 -220 11955
rect -290 11875 -275 11915
rect -235 11875 -220 11915
rect -290 11835 -220 11875
rect -290 11795 -275 11835
rect -235 11795 -220 11835
rect -290 11755 -220 11795
rect -290 11715 -275 11755
rect -235 11715 -220 11755
rect -290 11675 -220 11715
rect -290 11635 -275 11675
rect -235 11635 -220 11675
rect -290 11595 -220 11635
rect -290 11555 -275 11595
rect -235 11555 -220 11595
rect -290 11515 -220 11555
rect -290 11475 -275 11515
rect -235 11475 -220 11515
rect -290 11435 -220 11475
rect -290 11395 -275 11435
rect -235 11395 -220 11435
rect -290 11355 -220 11395
rect -290 11315 -275 11355
rect -235 11315 -220 11355
rect -290 11275 -220 11315
rect -290 11235 -275 11275
rect -235 11235 -220 11275
rect -290 11195 -220 11235
rect -290 11155 -275 11195
rect -235 11155 -220 11195
rect -290 11115 -220 11155
rect -290 11075 -275 11115
rect -235 11075 -220 11115
rect -290 11035 -220 11075
rect -290 10995 -275 11035
rect -235 10995 -220 11035
rect -290 10955 -220 10995
rect -290 10915 -275 10955
rect -235 10915 -220 10955
rect -290 10875 -220 10915
rect -290 10835 -275 10875
rect -235 10835 -220 10875
rect -290 10795 -220 10835
rect -290 10755 -275 10795
rect -235 10755 -220 10795
rect -290 10715 -220 10755
rect -290 10675 -275 10715
rect -235 10675 -220 10715
rect -290 10635 -220 10675
rect -290 10595 -275 10635
rect -235 10595 -220 10635
rect -290 10555 -220 10595
rect -290 10515 -275 10555
rect -235 10515 -220 10555
rect -290 10475 -220 10515
rect -290 10435 -275 10475
rect -235 10435 -220 10475
rect -290 10395 -220 10435
rect -290 10355 -275 10395
rect -235 10355 -220 10395
rect -290 10315 -220 10355
rect -290 10275 -275 10315
rect -235 10275 -220 10315
rect -290 10260 -220 10275
rect -345 10160 -305 10170
rect -345 10140 -335 10160
rect -315 10140 -305 10160
rect -345 10130 -305 10140
<< end >>
