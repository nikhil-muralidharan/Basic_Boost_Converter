magic
tech sky130A
timestamp 1640179460
<< nmos >>
rect -320 10245 -305 12270
<< ndiff >>
rect -420 12235 -320 12270
rect -420 12195 -390 12235
rect -350 12195 -320 12235
rect -420 12155 -320 12195
rect -420 12115 -390 12155
rect -350 12115 -320 12155
rect -420 12075 -320 12115
rect -420 12035 -390 12075
rect -350 12035 -320 12075
rect -420 11995 -320 12035
rect -420 11955 -390 11995
rect -350 11955 -320 11995
rect -420 11915 -320 11955
rect -420 11875 -390 11915
rect -350 11875 -320 11915
rect -420 11835 -320 11875
rect -420 11795 -390 11835
rect -350 11795 -320 11835
rect -420 11755 -320 11795
rect -420 11715 -390 11755
rect -350 11715 -320 11755
rect -420 11675 -320 11715
rect -420 11635 -390 11675
rect -350 11635 -320 11675
rect -420 11595 -320 11635
rect -420 11555 -390 11595
rect -350 11555 -320 11595
rect -420 11515 -320 11555
rect -420 11475 -390 11515
rect -350 11475 -320 11515
rect -420 11435 -320 11475
rect -420 11395 -390 11435
rect -350 11395 -320 11435
rect -420 11355 -320 11395
rect -420 11315 -390 11355
rect -350 11315 -320 11355
rect -420 11275 -320 11315
rect -420 11235 -390 11275
rect -350 11235 -320 11275
rect -420 11195 -320 11235
rect -420 11155 -390 11195
rect -350 11155 -320 11195
rect -420 11115 -320 11155
rect -420 11075 -390 11115
rect -350 11075 -320 11115
rect -420 11035 -320 11075
rect -420 10995 -390 11035
rect -350 10995 -320 11035
rect -420 10955 -320 10995
rect -420 10915 -390 10955
rect -350 10915 -320 10955
rect -420 10875 -320 10915
rect -420 10835 -390 10875
rect -350 10835 -320 10875
rect -420 10795 -320 10835
rect -420 10755 -390 10795
rect -350 10755 -320 10795
rect -420 10715 -320 10755
rect -420 10675 -390 10715
rect -350 10675 -320 10715
rect -420 10635 -320 10675
rect -420 10595 -390 10635
rect -350 10595 -320 10635
rect -420 10555 -320 10595
rect -420 10515 -390 10555
rect -350 10515 -320 10555
rect -420 10475 -320 10515
rect -420 10435 -390 10475
rect -350 10435 -320 10475
rect -420 10395 -320 10435
rect -420 10355 -390 10395
rect -350 10355 -320 10395
rect -420 10315 -320 10355
rect -420 10275 -390 10315
rect -350 10275 -320 10315
rect -420 10245 -320 10275
rect -305 12235 -205 12270
rect -305 12195 -275 12235
rect -235 12195 -205 12235
rect -305 12155 -205 12195
rect -305 12115 -275 12155
rect -235 12115 -205 12155
rect -305 12075 -205 12115
rect -305 12035 -275 12075
rect -235 12035 -205 12075
rect -305 11995 -205 12035
rect -305 11955 -275 11995
rect -235 11955 -205 11995
rect -305 11915 -205 11955
rect -305 11875 -275 11915
rect -235 11875 -205 11915
rect -305 11835 -205 11875
rect -305 11795 -275 11835
rect -235 11795 -205 11835
rect -305 11755 -205 11795
rect -305 11715 -275 11755
rect -235 11715 -205 11755
rect -305 11675 -205 11715
rect -305 11635 -275 11675
rect -235 11635 -205 11675
rect -305 11595 -205 11635
rect -305 11555 -275 11595
rect -235 11555 -205 11595
rect -305 11515 -205 11555
rect -305 11475 -275 11515
rect -235 11475 -205 11515
rect -305 11435 -205 11475
rect -305 11395 -275 11435
rect -235 11395 -205 11435
rect -305 11355 -205 11395
rect -305 11315 -275 11355
rect -235 11315 -205 11355
rect -305 11275 -205 11315
rect -305 11235 -275 11275
rect -235 11235 -205 11275
rect -305 11195 -205 11235
rect -305 11155 -275 11195
rect -235 11155 -205 11195
rect -305 11115 -205 11155
rect -305 11075 -275 11115
rect -235 11075 -205 11115
rect -305 11035 -205 11075
rect -305 10995 -275 11035
rect -235 10995 -205 11035
rect -305 10955 -205 10995
rect -305 10915 -275 10955
rect -235 10915 -205 10955
rect -305 10875 -205 10915
rect -305 10835 -275 10875
rect -235 10835 -205 10875
rect -305 10795 -205 10835
rect -305 10755 -275 10795
rect -235 10755 -205 10795
rect -305 10715 -205 10755
rect -305 10675 -275 10715
rect -235 10675 -205 10715
rect -305 10635 -205 10675
rect -305 10595 -275 10635
rect -235 10595 -205 10635
rect -305 10555 -205 10595
rect -305 10515 -275 10555
rect -235 10515 -205 10555
rect -305 10475 -205 10515
rect -305 10435 -275 10475
rect -235 10435 -205 10475
rect -305 10395 -205 10435
rect -305 10355 -275 10395
rect -235 10355 -205 10395
rect -305 10315 -205 10355
rect -305 10275 -275 10315
rect -235 10275 -205 10315
rect -305 10245 -205 10275
<< ndiffc >>
rect -390 12195 -350 12235
rect -390 12115 -350 12155
rect -390 12035 -350 12075
rect -390 11955 -350 11995
rect -390 11875 -350 11915
rect -390 11795 -350 11835
rect -390 11715 -350 11755
rect -390 11635 -350 11675
rect -390 11555 -350 11595
rect -390 11475 -350 11515
rect -390 11395 -350 11435
rect -390 11315 -350 11355
rect -390 11235 -350 11275
rect -390 11155 -350 11195
rect -390 11075 -350 11115
rect -390 10995 -350 11035
rect -390 10915 -350 10955
rect -390 10835 -350 10875
rect -390 10755 -350 10795
rect -390 10675 -350 10715
rect -390 10595 -350 10635
rect -390 10515 -350 10555
rect -390 10435 -350 10475
rect -390 10355 -350 10395
rect -390 10275 -350 10315
rect -275 12195 -235 12235
rect -275 12115 -235 12155
rect -275 12035 -235 12075
rect -275 11955 -235 11995
rect -275 11875 -235 11915
rect -275 11795 -235 11835
rect -275 11715 -235 11755
rect -275 11635 -235 11675
rect -275 11555 -235 11595
rect -275 11475 -235 11515
rect -275 11395 -235 11435
rect -275 11315 -235 11355
rect -275 11235 -235 11275
rect -275 11155 -235 11195
rect -275 11075 -235 11115
rect -275 10995 -235 11035
rect -275 10915 -235 10955
rect -275 10835 -235 10875
rect -275 10755 -235 10795
rect -275 10675 -235 10715
rect -275 10595 -235 10635
rect -275 10515 -235 10555
rect -275 10435 -235 10475
rect -275 10355 -235 10395
rect -275 10275 -235 10315
<< psubdiff >>
rect -520 12235 -420 12270
rect -520 12195 -490 12235
rect -450 12195 -420 12235
rect -520 12155 -420 12195
rect -520 12115 -490 12155
rect -450 12115 -420 12155
rect -520 12075 -420 12115
rect -520 12035 -490 12075
rect -450 12035 -420 12075
rect -520 11995 -420 12035
rect -520 11955 -490 11995
rect -450 11955 -420 11995
rect -520 11915 -420 11955
rect -520 11875 -490 11915
rect -450 11875 -420 11915
rect -520 11835 -420 11875
rect -520 11795 -490 11835
rect -450 11795 -420 11835
rect -520 11755 -420 11795
rect -520 11715 -490 11755
rect -450 11715 -420 11755
rect -520 11675 -420 11715
rect -520 11635 -490 11675
rect -450 11635 -420 11675
rect -520 11595 -420 11635
rect -520 11555 -490 11595
rect -450 11555 -420 11595
rect -520 11515 -420 11555
rect -520 11475 -490 11515
rect -450 11475 -420 11515
rect -520 11435 -420 11475
rect -520 11395 -490 11435
rect -450 11395 -420 11435
rect -520 11355 -420 11395
rect -520 11315 -490 11355
rect -450 11315 -420 11355
rect -520 11275 -420 11315
rect -520 11235 -490 11275
rect -450 11235 -420 11275
rect -520 11195 -420 11235
rect -520 11155 -490 11195
rect -450 11155 -420 11195
rect -520 11115 -420 11155
rect -520 11075 -490 11115
rect -450 11075 -420 11115
rect -520 11035 -420 11075
rect -520 10995 -490 11035
rect -450 10995 -420 11035
rect -520 10955 -420 10995
rect -520 10915 -490 10955
rect -450 10915 -420 10955
rect -520 10875 -420 10915
rect -520 10835 -490 10875
rect -450 10835 -420 10875
rect -520 10795 -420 10835
rect -520 10755 -490 10795
rect -450 10755 -420 10795
rect -520 10715 -420 10755
rect -520 10675 -490 10715
rect -450 10675 -420 10715
rect -520 10635 -420 10675
rect -520 10595 -490 10635
rect -450 10595 -420 10635
rect -520 10555 -420 10595
rect -520 10515 -490 10555
rect -450 10515 -420 10555
rect -520 10475 -420 10515
rect -520 10435 -490 10475
rect -450 10435 -420 10475
rect -520 10395 -420 10435
rect -520 10355 -490 10395
rect -450 10355 -420 10395
rect -520 10315 -420 10355
rect -520 10275 -490 10315
rect -450 10275 -420 10315
rect -520 10245 -420 10275
<< psubdiffcont >>
rect -490 12195 -450 12235
rect -490 12115 -450 12155
rect -490 12035 -450 12075
rect -490 11955 -450 11995
rect -490 11875 -450 11915
rect -490 11795 -450 11835
rect -490 11715 -450 11755
rect -490 11635 -450 11675
rect -490 11555 -450 11595
rect -490 11475 -450 11515
rect -490 11395 -450 11435
rect -490 11315 -450 11355
rect -490 11235 -450 11275
rect -490 11155 -450 11195
rect -490 11075 -450 11115
rect -490 10995 -450 11035
rect -490 10915 -450 10955
rect -490 10835 -450 10875
rect -490 10755 -450 10795
rect -490 10675 -450 10715
rect -490 10595 -450 10635
rect -490 10515 -450 10555
rect -490 10435 -450 10475
rect -490 10355 -450 10395
rect -490 10275 -450 10315
<< poly >>
rect -320 12270 -305 12290
rect -320 10170 -305 10245
rect -345 10160 -305 10170
rect -345 10140 -335 10160
rect -315 10140 -305 10160
rect -345 10130 -305 10140
<< polycont >>
rect -335 10140 -315 10160
<< locali >>
rect -505 12235 -335 12255
rect -505 12195 -490 12235
rect -450 12195 -390 12235
rect -350 12195 -335 12235
rect -505 12155 -335 12195
rect -505 12115 -490 12155
rect -450 12115 -390 12155
rect -350 12115 -335 12155
rect -505 12075 -335 12115
rect -505 12035 -490 12075
rect -450 12035 -390 12075
rect -350 12035 -335 12075
rect -505 11995 -335 12035
rect -505 11955 -490 11995
rect -450 11955 -390 11995
rect -350 11955 -335 11995
rect -505 11915 -335 11955
rect -505 11875 -490 11915
rect -450 11875 -390 11915
rect -350 11875 -335 11915
rect -505 11835 -335 11875
rect -505 11795 -490 11835
rect -450 11795 -390 11835
rect -350 11795 -335 11835
rect -505 11755 -335 11795
rect -505 11715 -490 11755
rect -450 11715 -390 11755
rect -350 11715 -335 11755
rect -505 11675 -335 11715
rect -505 11635 -490 11675
rect -450 11635 -390 11675
rect -350 11635 -335 11675
rect -505 11595 -335 11635
rect -505 11555 -490 11595
rect -450 11555 -390 11595
rect -350 11555 -335 11595
rect -505 11515 -335 11555
rect -505 11475 -490 11515
rect -450 11475 -390 11515
rect -350 11475 -335 11515
rect -505 11435 -335 11475
rect -505 11395 -490 11435
rect -450 11395 -390 11435
rect -350 11395 -335 11435
rect -505 11355 -335 11395
rect -505 11315 -490 11355
rect -450 11315 -390 11355
rect -350 11315 -335 11355
rect -505 11275 -335 11315
rect -505 11235 -490 11275
rect -450 11235 -390 11275
rect -350 11235 -335 11275
rect -505 11195 -335 11235
rect -505 11155 -490 11195
rect -450 11155 -390 11195
rect -350 11155 -335 11195
rect -505 11115 -335 11155
rect -505 11075 -490 11115
rect -450 11075 -390 11115
rect -350 11075 -335 11115
rect -505 11035 -335 11075
rect -505 10995 -490 11035
rect -450 10995 -390 11035
rect -350 10995 -335 11035
rect -505 10955 -335 10995
rect -505 10915 -490 10955
rect -450 10915 -390 10955
rect -350 10915 -335 10955
rect -505 10875 -335 10915
rect -505 10835 -490 10875
rect -450 10835 -390 10875
rect -350 10835 -335 10875
rect -505 10795 -335 10835
rect -505 10755 -490 10795
rect -450 10755 -390 10795
rect -350 10755 -335 10795
rect -505 10715 -335 10755
rect -505 10675 -490 10715
rect -450 10675 -390 10715
rect -350 10675 -335 10715
rect -505 10635 -335 10675
rect -505 10595 -490 10635
rect -450 10595 -390 10635
rect -350 10595 -335 10635
rect -505 10555 -335 10595
rect -505 10515 -490 10555
rect -450 10515 -390 10555
rect -350 10515 -335 10555
rect -505 10475 -335 10515
rect -505 10435 -490 10475
rect -450 10435 -390 10475
rect -350 10435 -335 10475
rect -505 10395 -335 10435
rect -505 10355 -490 10395
rect -450 10355 -390 10395
rect -350 10355 -335 10395
rect -505 10315 -335 10355
rect -505 10275 -490 10315
rect -450 10275 -390 10315
rect -350 10275 -335 10315
rect -505 10260 -335 10275
rect -290 12235 -220 12255
rect -290 12195 -275 12235
rect -235 12195 -220 12235
rect -290 12155 -220 12195
rect -290 12115 -275 12155
rect -235 12115 -220 12155
rect -290 12075 -220 12115
rect -290 12035 -275 12075
rect -235 12035 -220 12075
rect -290 11995 -220 12035
rect -290 11955 -275 11995
rect -235 11955 -220 11995
rect -290 11915 -220 11955
rect -290 11875 -275 11915
rect -235 11875 -220 11915
rect -290 11835 -220 11875
rect -290 11795 -275 11835
rect -235 11795 -220 11835
rect -290 11755 -220 11795
rect -290 11715 -275 11755
rect -235 11715 -220 11755
rect -290 11675 -220 11715
rect -290 11635 -275 11675
rect -235 11635 -220 11675
rect -290 11595 -220 11635
rect -290 11555 -275 11595
rect -235 11555 -220 11595
rect -290 11515 -220 11555
rect -290 11475 -275 11515
rect -235 11475 -220 11515
rect -290 11435 -220 11475
rect -290 11395 -275 11435
rect -235 11395 -220 11435
rect -290 11355 -220 11395
rect -290 11315 -275 11355
rect -235 11315 -220 11355
rect -290 11275 -220 11315
rect -290 11235 -275 11275
rect -235 11235 -220 11275
rect -290 11195 -220 11235
rect -290 11155 -275 11195
rect -235 11155 -220 11195
rect -290 11115 -220 11155
rect -290 11075 -275 11115
rect -235 11075 -220 11115
rect -290 11035 -220 11075
rect -290 10995 -275 11035
rect -235 10995 -220 11035
rect -290 10955 -220 10995
rect -290 10915 -275 10955
rect -235 10915 -220 10955
rect -290 10875 -220 10915
rect -290 10835 -275 10875
rect -235 10835 -220 10875
rect -290 10795 -220 10835
rect -290 10755 -275 10795
rect -235 10755 -220 10795
rect -290 10715 -220 10755
rect -290 10675 -275 10715
rect -235 10675 -220 10715
rect -290 10635 -220 10675
rect -290 10595 -275 10635
rect -235 10595 -220 10635
rect -290 10555 -220 10595
rect -290 10515 -275 10555
rect -235 10515 -220 10555
rect -290 10475 -220 10515
rect -290 10435 -275 10475
rect -235 10435 -220 10475
rect -290 10395 -220 10435
rect -290 10355 -275 10395
rect -235 10355 -220 10395
rect -290 10315 -220 10355
rect -290 10275 -275 10315
rect -235 10275 -220 10315
rect -290 10260 -220 10275
rect -345 10160 -305 10170
rect -345 10140 -335 10160
rect -315 10140 -305 10160
rect -345 10130 -305 10140
<< end >>
