magic
tech sky130A
timestamp 1659695591
<< nwell >>
rect -375 135 95 295
<< pmoslvt >>
rect -220 165 -185 265
rect -15 165 20 265
<< nmoslvt >>
rect -220 -120 -205 -20
rect -15 -120 0 -20
<< ndiff >>
rect -270 -35 -220 -20
rect -270 -105 -255 -35
rect -235 -105 -220 -35
rect -270 -120 -220 -105
rect -205 -35 -155 -20
rect -205 -105 -190 -35
rect -170 -105 -155 -35
rect -205 -120 -155 -105
rect -65 -35 -15 -20
rect -65 -105 -50 -35
rect -30 -105 -15 -35
rect -65 -120 -15 -105
rect 0 -35 50 -20
rect 0 -105 15 -35
rect 35 -105 50 -35
rect 0 -120 50 -105
<< pdiff >>
rect -270 250 -220 265
rect -270 180 -255 250
rect -235 180 -220 250
rect -270 165 -220 180
rect -185 250 -135 265
rect -185 180 -170 250
rect -150 180 -135 250
rect -185 165 -135 180
rect -65 250 -15 265
rect -65 180 -50 250
rect -30 180 -15 250
rect -65 165 -15 180
rect 20 250 70 265
rect 20 180 35 250
rect 55 180 70 250
rect 20 165 70 180
<< ndiffc >>
rect -255 -105 -235 -35
rect -190 -105 -170 -35
rect -50 -105 -30 -35
rect 15 -105 35 -35
<< pdiffc >>
rect -255 180 -235 250
rect -170 180 -150 250
rect -50 180 -30 250
rect 35 180 55 250
<< psubdiff >>
rect -355 -35 -305 -20
rect -355 -105 -340 -35
rect -320 -105 -305 -35
rect -355 -120 -305 -105
<< psubdiffcont >>
rect -340 -105 -320 -35
<< poly >>
rect -20 310 20 320
rect -20 290 -10 310
rect 10 290 20 310
rect -20 280 20 290
rect -220 265 -185 280
rect -15 265 20 280
rect -220 150 -185 165
rect -15 150 20 165
rect -240 140 -200 150
rect -240 120 -230 140
rect -210 120 -200 140
rect -240 110 -200 120
rect -245 25 -205 35
rect -245 5 -235 25
rect -215 5 -205 25
rect -245 -5 -205 5
rect -220 -20 -205 -5
rect -15 -20 0 -5
rect -220 -135 -205 -120
rect -15 -135 0 -120
rect -245 -145 -205 -135
rect -245 -165 -235 -145
rect -215 -165 -205 -145
rect -245 -175 -205 -165
rect -40 -145 0 -135
rect -40 -165 -30 -145
rect -10 -165 0 -145
rect -40 -175 0 -165
<< polycont >>
rect -10 290 10 310
rect -230 120 -210 140
rect -235 5 -215 25
rect -235 -165 -215 -145
rect -30 -165 -10 -145
<< locali >>
rect -20 310 20 320
rect -170 290 -10 310
rect 10 290 20 310
rect -170 260 -150 290
rect -20 280 20 290
rect -265 250 -225 260
rect -265 180 -255 250
rect -235 180 -225 250
rect -265 170 -225 180
rect -180 250 -140 260
rect -180 180 -170 250
rect -150 180 -140 250
rect -180 170 -140 180
rect -60 250 -20 260
rect -60 180 -50 250
rect -30 180 -20 250
rect -240 140 -200 150
rect -240 120 -230 140
rect -210 120 -200 140
rect -240 110 -200 120
rect -375 35 -335 45
rect -235 35 -210 110
rect -375 15 -365 35
rect -345 15 -335 35
rect -375 5 -335 15
rect -245 25 -205 35
rect -245 5 -235 25
rect -215 5 -205 25
rect -245 -5 -205 5
rect -180 -25 -160 170
rect -350 -35 -310 -25
rect -350 -105 -340 -35
rect -320 -105 -310 -35
rect -350 -115 -310 -105
rect -265 -35 -225 -25
rect -265 -105 -255 -35
rect -235 -105 -225 -35
rect -265 -115 -225 -105
rect -200 -35 -160 -25
rect -200 -105 -190 -35
rect -170 -105 -160 -35
rect -200 -115 -160 -105
rect -60 35 -20 180
rect 25 250 65 260
rect 25 180 35 250
rect 55 180 65 250
rect 25 170 65 180
rect 35 35 55 170
rect -60 15 -50 35
rect -30 15 -20 35
rect -60 -35 -20 15
rect 15 15 55 35
rect 15 -25 35 15
rect -60 -105 -50 -35
rect -30 -105 -20 -35
rect -60 -115 -20 -105
rect 5 -35 45 -25
rect 5 -105 15 -35
rect 35 -105 45 -35
rect 5 -115 45 -105
rect -375 -145 -205 -135
rect -40 -145 0 -135
rect -375 -155 -235 -145
rect -245 -165 -235 -155
rect -215 -165 -30 -145
rect -10 -165 0 -145
rect -245 -175 -205 -165
rect -40 -175 0 -165
rect 20 -175 40 -115
<< viali >>
rect -255 180 -235 250
rect -365 15 -345 35
rect -340 -105 -320 -35
rect -255 -105 -235 -35
rect -50 15 -30 35
<< metal1 >>
rect -375 250 95 260
rect -375 180 -255 250
rect -235 180 95 250
rect -375 170 95 180
rect -375 35 -20 45
rect -375 15 -365 35
rect -345 15 -50 35
rect -30 15 -20 35
rect -375 5 -20 15
rect -375 -35 95 -25
rect -375 -105 -340 -35
rect -320 -105 -255 -35
rect -235 -105 95 -35
rect -375 -115 95 -105
<< labels >>
rlabel metal1 -375 -70 -375 -70 7 VN
port 2 w
rlabel locali -375 -145 -375 -145 7 Control
port 3 w
rlabel metal1 -375 25 -375 25 7 Vin
port 4 w
rlabel metal1 -375 215 -375 215 7 VP
port 1 w
rlabel locali 30 -175 30 -175 5 Vout
port 5 s
<< end >>
