magic
tech sky130A
timestamp 1660234770
<< nwell >>
rect -280 95 490 240
<< nmos >>
rect -115 -75 -100 25
rect 55 -75 70 25
rect 225 -75 240 25
rect 395 -75 410 25
<< pmoslvt >>
rect -125 120 -90 220
rect 45 120 80 220
rect 215 120 250 220
rect 385 120 420 220
<< ndiff >>
rect -165 10 -115 25
rect -165 -60 -150 10
rect -130 -60 -115 10
rect -165 -75 -115 -60
rect -100 10 55 25
rect -100 -60 -85 10
rect -65 -60 20 10
rect 40 -60 55 10
rect -100 -75 55 -60
rect 70 10 225 25
rect 70 -60 85 10
rect 105 -60 190 10
rect 210 -60 225 10
rect 70 -75 225 -60
rect 240 10 395 25
rect 240 -60 255 10
rect 275 -60 360 10
rect 380 -60 395 10
rect 240 -75 395 -60
rect 410 10 460 25
rect 410 -60 425 10
rect 445 -60 460 10
rect 410 -75 460 -60
<< pdiff >>
rect -175 205 -125 220
rect -175 135 -160 205
rect -140 135 -125 205
rect -175 120 -125 135
rect -90 205 -40 220
rect -90 135 -75 205
rect -55 135 -40 205
rect -90 120 -40 135
rect -5 205 45 220
rect -5 135 10 205
rect 30 135 45 205
rect -5 120 45 135
rect 80 205 130 220
rect 80 135 95 205
rect 115 135 130 205
rect 80 120 130 135
rect 165 205 215 220
rect 165 135 180 205
rect 200 135 215 205
rect 165 120 215 135
rect 250 205 300 220
rect 250 135 265 205
rect 285 135 300 205
rect 250 120 300 135
rect 335 205 385 220
rect 335 135 350 205
rect 370 135 385 205
rect 335 120 385 135
rect 420 205 470 220
rect 420 135 435 205
rect 455 135 470 205
rect 420 120 470 135
<< ndiffc >>
rect -150 -60 -130 10
rect -85 -60 -65 10
rect 20 -60 40 10
rect 85 -60 105 10
rect 190 -60 210 10
rect 255 -60 275 10
rect 360 -60 380 10
rect 425 -60 445 10
<< pdiffc >>
rect -160 135 -140 205
rect -75 135 -55 205
rect 10 135 30 205
rect 95 135 115 205
rect 180 135 200 205
rect 265 135 285 205
rect 350 135 370 205
rect 435 135 455 205
<< psubdiff >>
rect -255 10 -205 25
rect -255 -60 -240 10
rect -220 -60 -205 10
rect -255 -75 -205 -60
<< nsubdiff >>
rect -260 205 -210 220
rect -260 135 -245 205
rect -225 135 -210 205
rect -260 120 -210 135
<< psubdiffcont >>
rect -240 -60 -220 10
<< nsubdiffcont >>
rect -245 135 -225 205
<< poly >>
rect -125 220 -90 235
rect 45 220 80 235
rect 215 220 250 235
rect 385 220 420 235
rect -125 105 -90 120
rect 45 105 80 120
rect 215 105 250 120
rect 385 105 420 120
rect -115 25 -100 105
rect 55 80 70 105
rect 225 80 240 105
rect 55 70 95 80
rect 55 50 65 70
rect 85 50 95 70
rect 55 40 95 50
rect 200 70 240 80
rect 200 50 210 70
rect 230 50 240 70
rect 200 40 240 50
rect 55 25 70 40
rect 225 25 240 40
rect 395 25 410 105
rect -115 -90 -100 -75
rect 55 -90 70 -75
rect 225 -90 240 -75
rect 395 -90 410 -75
rect -140 -100 -100 -90
rect -140 -120 -130 -100
rect -110 -120 -100 -100
rect -140 -130 -100 -120
rect 30 -100 70 -90
rect 30 -120 40 -100
rect 60 -120 70 -100
rect 30 -130 70 -120
rect 200 -100 240 -90
rect 200 -120 210 -100
rect 230 -120 240 -100
rect 200 -130 240 -120
rect 370 -100 410 -90
rect 370 -120 380 -100
rect 400 -120 410 -100
rect 370 -130 410 -120
<< polycont >>
rect 65 50 85 70
rect 210 50 230 70
rect -130 -120 -110 -100
rect 40 -120 60 -100
rect 210 -120 230 -100
rect 380 -120 400 -100
<< locali >>
rect -255 205 -215 215
rect -255 135 -245 205
rect -225 135 -215 205
rect -255 125 -215 135
rect -170 205 -130 215
rect -170 135 -160 205
rect -140 135 -130 205
rect -170 125 -130 135
rect -85 205 -45 215
rect -85 135 -75 205
rect -55 135 -45 205
rect -85 125 -45 135
rect 0 205 40 215
rect 0 135 10 205
rect 30 135 40 205
rect 0 125 40 135
rect 85 205 125 215
rect 85 135 95 205
rect 115 135 125 205
rect 85 125 125 135
rect 170 205 210 215
rect 170 135 180 205
rect 200 135 210 205
rect 170 125 210 135
rect 255 205 295 215
rect 255 135 265 205
rect 285 135 295 205
rect 255 125 295 135
rect 340 205 380 215
rect 340 135 350 205
rect 370 135 380 205
rect 340 125 380 135
rect 425 205 465 215
rect 425 135 435 205
rect 455 135 465 205
rect 425 125 465 135
rect -75 90 -55 125
rect 10 90 30 125
rect 265 90 285 125
rect 435 90 455 125
rect -75 70 105 90
rect 55 50 65 70
rect 85 50 105 70
rect 55 40 105 50
rect 85 20 105 40
rect 190 70 455 90
rect 190 50 210 70
rect 230 50 240 70
rect 190 40 240 50
rect 190 20 210 40
rect -250 10 -210 20
rect -250 -60 -240 10
rect -220 -60 -210 10
rect -250 -70 -210 -60
rect -160 10 -120 20
rect -160 -60 -150 10
rect -130 -60 -120 10
rect -160 -70 -120 -60
rect -95 10 50 20
rect -95 -60 -85 10
rect -65 -60 20 10
rect 40 -60 50 10
rect -95 -65 50 -60
rect 75 10 115 20
rect 75 -60 85 10
rect 105 -60 115 10
rect 75 -65 115 -60
rect 180 10 220 20
rect 180 -60 190 10
rect 210 -60 220 10
rect 180 -65 220 -60
rect 245 10 390 20
rect 245 -60 255 10
rect 275 -60 360 10
rect 380 -60 390 10
rect 245 -65 390 -60
rect 415 10 455 20
rect 415 -60 425 10
rect 445 -60 455 10
rect 415 -65 455 -60
rect -140 -100 -100 -90
rect -140 -120 -130 -100
rect -110 -120 -100 -100
rect -140 -130 -100 -120
rect 30 -100 70 -90
rect 30 -120 40 -100
rect 60 -120 70 -100
rect 30 -130 70 -120
rect 200 -100 240 -90
rect 200 -120 210 -100
rect 230 -120 240 -100
rect 200 -130 240 -120
rect 370 -100 410 -90
rect 370 -120 380 -100
rect 400 -120 410 -100
rect 370 -130 410 -120
<< viali >>
rect -245 135 -225 205
rect -75 135 -55 205
rect 95 135 115 205
rect 180 135 200 205
rect 350 135 370 205
rect -150 -60 -130 10
rect 425 -60 445 10
<< metal1 >>
rect -280 205 490 215
rect -280 135 -245 205
rect -225 135 -75 205
rect -55 135 95 205
rect 115 135 180 205
rect 200 135 350 205
rect 370 135 490 205
rect -280 125 490 135
rect -280 10 500 20
rect -280 -60 -150 10
rect -130 -60 425 10
rect 445 -60 500 10
rect -280 -70 500 -60
<< labels >>
rlabel metal1 -280 170 -280 170 7 VP
port 1 w
rlabel metal1 -280 -20 -280 -20 7 VN
port 2 w
rlabel locali -120 -130 -120 -130 5 S
port 3 s
rlabel locali 50 -130 50 -130 5 Q
port 5 s
rlabel locali 220 -130 220 -130 5 Qb
port 6 s
rlabel locali 390 -130 390 -130 5 R
port 4 s
<< end >>
