magic
tech sky130A
timestamp 1660760052
<< nwell >>
rect -280 95 490 240
<< nmos >>
rect -115 -350 -100 -250
rect 55 -350 70 -250
rect 225 -350 240 -250
rect 395 -350 410 -250
<< pmoslvt >>
rect -125 120 -90 220
rect 45 120 80 220
rect 215 120 250 220
rect 385 120 420 220
<< ndiff >>
rect -165 -265 -115 -250
rect -165 -335 -150 -265
rect -130 -335 -115 -265
rect -165 -350 -115 -335
rect -100 -265 55 -250
rect -100 -335 -85 -265
rect -65 -335 20 -265
rect 40 -335 55 -265
rect -100 -350 55 -335
rect 70 -265 225 -250
rect 70 -335 85 -265
rect 105 -335 190 -265
rect 210 -335 225 -265
rect 70 -350 225 -335
rect 240 -265 395 -250
rect 240 -335 255 -265
rect 275 -335 360 -265
rect 380 -335 395 -265
rect 240 -350 395 -335
rect 410 -265 460 -250
rect 410 -335 425 -265
rect 445 -335 460 -265
rect 410 -350 460 -335
<< pdiff >>
rect -175 205 -125 220
rect -175 135 -160 205
rect -140 135 -125 205
rect -175 120 -125 135
rect -90 205 -40 220
rect -90 135 -75 205
rect -55 135 -40 205
rect -90 120 -40 135
rect -5 205 45 220
rect -5 135 10 205
rect 30 135 45 205
rect -5 120 45 135
rect 80 205 130 220
rect 80 135 95 205
rect 115 135 130 205
rect 80 120 130 135
rect 165 205 215 220
rect 165 135 180 205
rect 200 135 215 205
rect 165 120 215 135
rect 250 205 300 220
rect 250 135 265 205
rect 285 135 300 205
rect 250 120 300 135
rect 335 205 385 220
rect 335 135 350 205
rect 370 135 385 205
rect 335 120 385 135
rect 420 205 470 220
rect 420 135 435 205
rect 455 135 470 205
rect 420 120 470 135
<< ndiffc >>
rect -150 -335 -130 -265
rect -85 -335 -65 -265
rect 20 -335 40 -265
rect 85 -335 105 -265
rect 190 -335 210 -265
rect 255 -335 275 -265
rect 360 -335 380 -265
rect 425 -335 445 -265
<< pdiffc >>
rect -160 135 -140 205
rect -75 135 -55 205
rect 10 135 30 205
rect 95 135 115 205
rect 180 135 200 205
rect 265 135 285 205
rect 350 135 370 205
rect 435 135 455 205
<< psubdiff >>
rect -255 -265 -205 -250
rect -255 -335 -240 -265
rect -220 -335 -205 -265
rect -255 -350 -205 -335
<< nsubdiff >>
rect -260 205 -210 220
rect -260 135 -245 205
rect -225 135 -210 205
rect -260 120 -210 135
<< psubdiffcont >>
rect -240 -335 -220 -265
<< nsubdiffcont >>
rect -245 135 -225 205
<< poly >>
rect -125 220 -90 235
rect 45 220 80 235
rect 215 220 250 235
rect 385 220 420 235
rect -125 105 -90 120
rect 45 105 80 120
rect 215 105 250 120
rect 385 105 420 120
rect -115 25 -100 105
rect 55 80 70 105
rect 225 80 240 105
rect 55 70 95 80
rect 55 50 65 70
rect 85 50 95 70
rect 55 40 95 50
rect 200 70 240 80
rect 200 50 210 70
rect 230 50 240 70
rect 200 40 240 50
rect -140 15 -100 25
rect -140 -5 -130 15
rect -110 -5 -100 15
rect -140 -15 -100 -5
rect 395 25 410 105
rect 395 15 435 25
rect 395 -5 405 15
rect 425 -5 435 15
rect 395 -15 435 -5
rect -140 -205 -100 -195
rect -140 -225 -130 -205
rect -110 -225 -100 -205
rect -140 -235 -100 -225
rect -115 -250 -100 -235
rect 55 -205 95 -195
rect 55 -225 65 -205
rect 85 -225 95 -205
rect 55 -235 95 -225
rect 200 -205 240 -195
rect 200 -225 210 -205
rect 230 -225 240 -205
rect 200 -235 240 -225
rect 55 -250 70 -235
rect 225 -250 240 -235
rect 395 -205 435 -195
rect 395 -225 405 -205
rect 425 -225 435 -205
rect 395 -235 435 -225
rect 395 -250 410 -235
rect -115 -365 -100 -350
rect 55 -365 70 -350
rect 225 -365 240 -350
rect 395 -365 410 -350
rect -140 -375 -100 -365
rect -140 -395 -130 -375
rect -110 -395 -100 -375
rect -140 -405 -100 -395
rect 30 -375 70 -365
rect 30 -395 40 -375
rect 60 -395 70 -375
rect 30 -405 70 -395
rect 200 -375 240 -365
rect 200 -395 210 -375
rect 230 -395 240 -375
rect 200 -405 240 -395
rect 370 -375 410 -365
rect 370 -395 380 -375
rect 400 -395 410 -375
rect 370 -405 410 -395
<< polycont >>
rect 65 50 85 70
rect 210 50 230 70
rect -130 -5 -110 15
rect 405 -5 425 15
rect -130 -225 -110 -205
rect 65 -225 85 -205
rect 210 -225 230 -205
rect 405 -225 425 -205
rect -130 -395 -110 -375
rect 40 -395 60 -375
rect 210 -395 230 -375
rect 380 -395 400 -375
<< locali >>
rect -255 205 -215 215
rect -255 135 -245 205
rect -225 135 -215 205
rect -255 125 -215 135
rect -170 205 -130 215
rect -170 135 -160 205
rect -140 135 -130 205
rect -170 125 -130 135
rect -85 205 -45 215
rect -85 135 -75 205
rect -55 135 -45 205
rect -85 125 -45 135
rect 0 205 40 215
rect 0 135 10 205
rect 30 135 40 205
rect 0 125 40 135
rect 85 205 125 215
rect 85 135 95 205
rect 115 135 125 205
rect 85 125 125 135
rect 170 205 210 215
rect 170 135 180 205
rect 200 135 210 205
rect 170 125 210 135
rect 255 205 295 215
rect 255 135 265 205
rect 285 135 295 205
rect 255 125 295 135
rect 340 205 380 215
rect 340 135 350 205
rect 370 135 380 205
rect 340 125 380 135
rect 425 205 465 215
rect 425 135 435 205
rect 455 135 465 205
rect 425 125 465 135
rect -75 90 -55 125
rect 10 90 30 125
rect 265 90 285 125
rect 435 90 455 125
rect -75 70 105 90
rect 55 50 65 70
rect 85 50 105 70
rect 55 40 105 50
rect -140 15 -100 25
rect -140 -5 -130 15
rect -110 -5 -100 15
rect -140 -15 -100 -5
rect -130 -195 -110 -15
rect 85 -195 105 40
rect -140 -205 -100 -195
rect -140 -225 -130 -205
rect -110 -225 -100 -205
rect -140 -235 -100 -225
rect 55 -205 105 -195
rect 55 -225 65 -205
rect 85 -225 105 -205
rect 55 -235 105 -225
rect 85 -255 105 -235
rect 190 70 455 90
rect 190 50 210 70
rect 230 50 240 70
rect 190 40 240 50
rect 190 -195 210 40
rect 395 15 435 25
rect 395 -5 405 15
rect 425 -5 435 15
rect 395 -15 435 -5
rect 405 -195 425 -15
rect 190 -205 240 -195
rect 190 -225 210 -205
rect 230 -225 240 -205
rect 190 -235 240 -225
rect 395 -205 435 -195
rect 395 -225 405 -205
rect 425 -225 435 -205
rect 395 -235 435 -225
rect 190 -255 210 -235
rect -250 -265 -210 -255
rect -250 -335 -240 -265
rect -220 -335 -210 -265
rect -250 -345 -210 -335
rect -160 -265 -120 -255
rect -160 -335 -150 -265
rect -130 -335 -120 -265
rect -160 -345 -120 -335
rect -95 -265 50 -255
rect -95 -335 -85 -265
rect -65 -335 20 -265
rect 40 -335 50 -265
rect -95 -340 50 -335
rect 75 -265 115 -255
rect 75 -335 85 -265
rect 105 -335 115 -265
rect 75 -340 115 -335
rect 180 -265 220 -255
rect 180 -335 190 -265
rect 210 -335 220 -265
rect 180 -340 220 -335
rect 245 -265 390 -255
rect 245 -335 255 -265
rect 275 -335 360 -265
rect 380 -335 390 -265
rect 245 -340 390 -335
rect 415 -265 455 -255
rect 415 -335 425 -265
rect 445 -335 455 -265
rect 415 -340 455 -335
rect -140 -375 -100 -365
rect -140 -395 -130 -375
rect -110 -395 -100 -375
rect -140 -405 -100 -395
rect 30 -375 70 -365
rect 30 -395 40 -375
rect 60 -395 70 -375
rect 30 -405 70 -395
rect 200 -375 240 -365
rect 200 -395 210 -375
rect 230 -395 240 -375
rect 200 -405 240 -395
rect 370 -375 410 -365
rect 370 -395 380 -375
rect 400 -395 410 -375
rect 370 -405 410 -395
<< viali >>
rect -245 135 -225 205
rect -75 135 -55 205
rect 95 135 115 205
rect 180 135 200 205
rect 350 135 370 205
rect -150 -335 -130 -265
rect 425 -335 445 -265
<< metal1 >>
rect -280 205 490 215
rect -280 135 -245 205
rect -225 135 -75 205
rect -55 135 95 205
rect 115 135 180 205
rect 200 135 350 205
rect 370 135 490 205
rect -280 125 490 135
rect -280 -265 505 -255
rect -280 -335 -150 -265
rect -130 -335 425 -265
rect 445 -335 505 -265
rect -280 -345 505 -335
<< labels >>
rlabel metal1 -280 170 -280 170 7 VP
port 1 w
rlabel metal1 -280 -295 -280 -295 7 VN
port 2 w
rlabel locali -120 -405 -120 -405 5 S
port 3 s
rlabel locali 50 -405 50 -405 5 Q
port 5 s
rlabel locali 220 -405 220 -405 5 Qb
port 6 s
rlabel locali 390 -405 390 -405 5 R
port 4 s
<< end >>
