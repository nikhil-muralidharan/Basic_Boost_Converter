magic
tech sky130A
timestamp 1657335720
<< nwell >>
rect -320 95 180 265
<< pmoslvt >>
rect -140 115 -105 245
rect 50 115 85 245
<< nmoslvt >>
rect -125 -45 -105 60
rect 70 -45 90 60
<< ndiff >>
rect -185 45 -125 60
rect -185 -25 -165 45
rect -140 -25 -125 45
rect -185 -45 -125 -25
rect -105 45 -45 60
rect -105 -25 -85 45
rect -60 -25 -45 45
rect -105 -45 -45 -25
rect 5 45 70 60
rect 5 -25 25 45
rect 50 -25 70 45
rect 5 -45 70 -25
rect 90 45 145 60
rect 90 -25 105 45
rect 130 -25 145 45
rect 90 -45 145 -25
<< pdiff >>
rect -185 230 -140 245
rect -185 135 -175 230
rect -150 135 -140 230
rect -185 115 -140 135
rect -105 230 -55 245
rect -105 135 -90 230
rect -65 135 -55 230
rect -105 115 -55 135
rect 5 230 50 245
rect 5 135 15 230
rect 40 135 50 230
rect 5 115 50 135
rect 85 230 135 245
rect 85 135 100 230
rect 125 135 135 230
rect 85 115 135 135
<< ndiffc >>
rect -165 -25 -140 45
rect -85 -25 -60 45
rect 25 -25 50 45
rect 105 -25 130 45
<< pdiffc >>
rect -175 135 -150 230
rect -90 135 -65 230
rect 15 135 40 230
rect 100 135 125 230
<< psubdiff >>
rect -295 45 -220 60
rect -295 -30 -270 45
rect -240 -30 -220 45
rect -295 -45 -220 -30
<< nsubdiff >>
rect -295 230 -220 245
rect -295 135 -270 230
rect -240 135 -220 230
rect -295 115 -220 135
<< psubdiffcont >>
rect -270 -30 -240 45
<< nsubdiffcont >>
rect -270 135 -240 230
<< poly >>
rect -140 245 -105 260
rect 50 245 85 260
rect -140 100 -105 115
rect -125 60 -105 100
rect 50 95 85 115
rect 70 60 90 95
rect -125 -60 -105 -45
rect 70 -60 90 -45
rect -125 -70 -85 -60
rect -125 -90 -115 -70
rect -95 -90 -85 -70
rect -125 -100 -85 -90
rect 70 -70 110 -60
rect 70 -90 80 -70
rect 100 -90 110 -70
rect 70 -100 110 -90
<< polycont >>
rect -115 -90 -95 -70
rect 80 -90 100 -70
<< locali >>
rect -280 230 -230 240
rect -280 135 -270 230
rect -240 135 -230 230
rect -280 125 -230 135
rect -180 230 -145 240
rect -180 135 -175 230
rect -150 135 -145 230
rect -180 125 -145 135
rect -95 230 -60 240
rect -95 135 -90 230
rect -65 135 -60 230
rect -95 100 -60 135
rect 10 230 45 240
rect 10 135 15 230
rect 40 135 45 230
rect 10 125 45 135
rect 95 230 130 240
rect 95 135 100 230
rect 125 135 130 230
rect 95 100 130 135
rect -95 75 180 100
rect -285 45 -230 55
rect -285 -30 -270 45
rect -240 -30 -230 45
rect -285 -40 -230 -30
rect -185 45 -130 55
rect -185 -25 -165 45
rect -140 -25 -130 45
rect -185 -35 -130 -25
rect -95 45 -50 75
rect -95 -25 -85 45
rect -60 -25 -50 45
rect -95 -35 -50 -25
rect 15 45 60 55
rect 15 -25 25 45
rect 50 -25 60 45
rect 15 -35 60 -25
rect 95 45 140 75
rect 95 -25 105 45
rect 130 -25 140 45
rect 95 -35 140 -25
rect -125 -70 -85 -60
rect -125 -90 -115 -70
rect -95 -90 -85 -70
rect -125 -100 -85 -90
rect 70 -70 110 -60
rect 70 -90 80 -70
rect 100 -90 110 -70
rect 70 -100 110 -90
<< viali >>
rect -270 135 -240 230
rect -175 135 -150 230
rect 15 135 40 230
rect -270 -30 -240 45
rect -165 -25 -140 45
rect 25 -25 50 45
<< metal1 >>
rect -320 230 180 240
rect -320 135 -270 230
rect -240 135 -175 230
rect -150 135 15 230
rect 40 135 180 230
rect -320 120 180 135
rect -320 45 180 55
rect -320 -30 -270 45
rect -240 -25 -165 45
rect -140 -25 25 45
rect 50 -25 180 45
rect -240 -30 180 -25
rect -320 -40 180 -30
<< labels >>
rlabel poly -120 70 -120 70 7 A
rlabel poly 80 65 80 65 7 B
rlabel metal1 -320 175 -320 175 7 VDD
rlabel metal1 -320 0 -320 0 7 GND
rlabel locali 180 90 180 90 7 Y
<< end >>
