magic
tech sky130A
timestamp 1659603320
<< nwell >>
rect -375 45 95 205
<< pmoslvt >>
rect -220 75 -185 175
rect -15 75 20 175
<< nmoslvt >>
rect -220 -120 -205 -20
rect -15 -120 0 -20
<< ndiff >>
rect -270 -35 -220 -20
rect -270 -105 -255 -35
rect -235 -105 -220 -35
rect -270 -120 -220 -105
rect -205 -35 -155 -20
rect -205 -105 -190 -35
rect -170 -105 -155 -35
rect -205 -120 -155 -105
rect -65 -35 -15 -20
rect -65 -105 -50 -35
rect -30 -105 -15 -35
rect -65 -120 -15 -105
rect 0 -35 50 -20
rect 0 -105 15 -35
rect 35 -105 50 -35
rect 0 -120 50 -105
<< pdiff >>
rect -270 160 -220 175
rect -270 90 -255 160
rect -235 90 -220 160
rect -270 75 -220 90
rect -185 160 -135 175
rect -185 90 -170 160
rect -150 90 -135 160
rect -185 75 -135 90
rect -65 160 -15 175
rect -65 90 -50 160
rect -30 90 -15 160
rect -65 75 -15 90
rect 20 160 70 175
rect 20 90 35 160
rect 55 90 70 160
rect 20 75 70 90
<< ndiffc >>
rect -255 -105 -235 -35
rect -190 -105 -170 -35
rect -50 -105 -30 -35
rect 15 -105 35 -35
<< pdiffc >>
rect -255 90 -235 160
rect -170 90 -150 160
rect -50 90 -30 160
rect 35 90 55 160
<< psubdiff >>
rect -355 -35 -305 -20
rect -355 -105 -340 -35
rect -320 -105 -305 -35
rect -355 -120 -305 -105
<< nsubdiff >>
rect -355 160 -305 175
rect -355 90 -340 160
rect -320 90 -305 160
rect -355 75 -305 90
<< psubdiffcont >>
rect -340 -105 -320 -35
<< nsubdiffcont >>
rect -340 90 -320 160
<< poly >>
rect -20 220 20 230
rect -20 200 -10 220
rect 10 200 20 220
rect -20 190 20 200
rect -220 175 -185 190
rect -15 175 20 190
rect -220 60 -185 75
rect -15 60 20 75
rect -220 -20 -205 60
rect -15 -20 0 -5
rect -220 -135 -205 -120
rect -15 -135 0 -120
rect -245 -145 -205 -135
rect -245 -165 -235 -145
rect -215 -165 -205 -145
rect -245 -175 -205 -165
rect -40 -145 0 -135
rect -40 -165 -30 -145
rect -10 -165 0 -145
rect -40 -175 0 -165
<< polycont >>
rect -10 200 10 220
rect -235 -165 -215 -145
rect -30 -165 -10 -145
<< locali >>
rect -20 220 20 230
rect -170 200 -10 220
rect 10 200 20 220
rect -170 170 -150 200
rect -20 190 20 200
rect -350 160 -310 170
rect -350 90 -340 160
rect -320 90 -310 160
rect -350 80 -310 90
rect -265 160 -225 170
rect -265 90 -255 160
rect -235 90 -225 160
rect -265 80 -225 90
rect -180 160 -140 170
rect -180 90 -170 160
rect -150 90 -140 160
rect -180 80 -140 90
rect -60 160 -20 170
rect -60 90 -50 160
rect -30 90 -20 160
rect -375 35 -335 45
rect -375 15 -365 35
rect -345 15 -335 35
rect -375 5 -335 15
rect -180 -25 -160 80
rect -350 -35 -310 -25
rect -350 -105 -340 -35
rect -320 -105 -310 -35
rect -350 -115 -310 -105
rect -265 -35 -225 -25
rect -265 -105 -255 -35
rect -235 -105 -225 -35
rect -265 -115 -225 -105
rect -200 -35 -160 -25
rect -200 -105 -190 -35
rect -170 -105 -160 -35
rect -200 -115 -160 -105
rect -60 35 -20 90
rect 25 160 65 170
rect 25 90 35 160
rect 55 90 65 160
rect 25 80 65 90
rect 35 35 55 80
rect -60 15 -50 35
rect -30 15 -20 35
rect -60 -35 -20 15
rect 15 15 95 35
rect 15 -25 35 15
rect -60 -105 -50 -35
rect -30 -105 -20 -35
rect -60 -115 -20 -105
rect 5 -35 45 -25
rect 5 -105 15 -35
rect 35 -105 45 -35
rect 5 -115 45 -105
rect -375 -145 -205 -135
rect -40 -145 0 -135
rect -375 -155 -235 -145
rect -245 -165 -235 -155
rect -215 -165 -30 -145
rect -10 -165 0 -145
rect -245 -175 -205 -165
rect -40 -175 0 -165
<< viali >>
rect -340 90 -320 160
rect -255 90 -235 160
rect -365 15 -345 35
rect -340 -105 -320 -35
rect -255 -105 -235 -35
rect -50 15 -30 35
<< metal1 >>
rect -375 160 95 170
rect -375 90 -340 160
rect -320 90 -255 160
rect -235 90 95 160
rect -375 80 95 90
rect -375 35 -20 45
rect -375 15 -365 35
rect -345 15 -50 35
rect -30 15 -20 35
rect -375 5 -20 15
rect -375 -35 95 -25
rect -375 -105 -340 -35
rect -320 -105 -255 -35
rect -235 -105 95 -35
rect -375 -115 95 -105
<< labels >>
rlabel metal1 -375 125 -375 125 7 VP
port 1 w
rlabel metal1 -375 -70 -375 -70 7 VN
port 2 w
rlabel locali -375 -145 -375 -145 7 Control
port 3 w
rlabel metal1 -375 25 -375 25 7 Vin
port 4 w
rlabel locali 95 25 95 25 3 Vout
port 5 e
<< end >>
